
module s38417 ( CK, g1249, g16297, g16355, g16399, g16437, g16496, g1943, 
        g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g2637, 
        g27380, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, 
        g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, 
        g3231, g3232, g3233, g3234, g3993, g4088, g4090, g4200, g4321, g4323, 
        g4450, g4590, g51, g5388, g5437, g5472, g5511, g5549, g5555, g5595, 
        g5612, g5629, g563, g5637, g5648, g5657, g5686, g5695, g5738, g5747, 
        g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, 
        g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, 
        g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, 
        g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, 
        g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, 
        g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, 
        g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, test_se, 
        test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, 
        test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, 
        test_si8, test_so8, test_si9, test_so9, test_si10, test_so10, 
        test_si11, test_so11, test_si12, test_so12, test_si13, test_so13, 
        test_si14, test_so14, test_si15, test_so15, test_si16, test_so16, 
        test_si17, test_so17, test_si18, test_so18, test_si19, test_so19, 
        test_si20, test_so20, test_si21, test_so21, test_si22, test_so22, 
        test_si23, test_so23, test_si24, test_so24, test_si25, test_so25, 
        test_si26, test_so26, test_si27, test_so27, test_si28, test_so28, 
        test_si29, test_so29, test_si30, test_so30, test_si31, test_so31, 
        test_si32, test_so32, test_si33, test_so33, test_si34, test_so34, 
        test_si35, test_so35, test_si36, test_so36, test_si37, test_so37, 
        test_si38, test_so38, test_si39, test_so39, test_si40, test_so40, 
        test_si41, test_so41, test_si42, test_so42, test_si43, test_so43, 
        test_si44, test_so44, test_si45, test_so45, test_si46, test_so46, 
        test_si47, test_so47, test_si48, test_so48, test_si49, test_so49, 
        test_si50, test_so50, test_si51, test_so51, test_si52, test_so52, 
        test_si53, test_so53, test_si54, test_so54, test_si55, test_so55, 
        test_si56, test_so56, test_si57, test_so57, test_si58, test_so58, 
        test_si59, test_so59, test_si60, test_so60, test_si61, test_so61, 
        test_si62, test_so62, test_si63, test_so63, test_si64, test_so64, 
        test_si65, test_so65, test_si66, test_so66, test_si67, test_so67, 
        test_si68, test_so68, test_si69, test_so69, test_si70, test_so70, 
        test_si71, test_so71, test_si72, test_so72, test_si73, test_so73, 
        test_si74, test_so74, test_si75, test_so75, test_si76, test_so76, 
        test_si77, test_so77, test_si78, test_so78, test_si79, test_so79, 
        test_si80, test_so80, test_si81, test_so81, test_si82, test_so82, 
        test_si83, test_so83, test_si84, test_so84, test_si85, test_so85, 
        test_si86, test_so86, test_si87, test_so87, test_si88, test_so88, 
        test_si89, test_so89, test_si90, test_so90, test_si91, test_so91, 
        test_si92, test_so92, test_si93, test_so93, test_si94, test_so94, 
        test_si95, test_so95, test_si96, test_so96, test_si97, test_so97, 
        test_si98, test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217,
         g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227,
         g3228, g3229, g3230, g3231, g3232, g3233, g3234, g51, g563, test_se,
         test_si1, test_si2, test_si3, test_si4, test_si5, test_si6, test_si7,
         test_si8, test_si9, test_si10, test_si11, test_si12, test_si13,
         test_si14, test_si15, test_si16, test_si17, test_si18, test_si19,
         test_si20, test_si21, test_si22, test_si23, test_si24, test_si25,
         test_si26, test_si27, test_si28, test_si29, test_si30, test_si31,
         test_si32, test_si33, test_si34, test_si35, test_si36, test_si37,
         test_si38, test_si39, test_si40, test_si41, test_si42, test_si43,
         test_si44, test_si45, test_si46, test_si47, test_si48, test_si49,
         test_si50, test_si51, test_si52, test_si53, test_si54, test_si55,
         test_si56, test_si57, test_si58, test_si59, test_si60, test_si61,
         test_si62, test_si63, test_si64, test_si65, test_si66, test_si67,
         test_si68, test_si69, test_si70, test_si71, test_si72, test_si73,
         test_si74, test_si75, test_si76, test_si77, test_si78, test_si79,
         test_si80, test_si81, test_si82, test_si83, test_si84, test_si85,
         test_si86, test_si87, test_si88, test_si89, test_si90, test_si91,
         test_si92, test_si93, test_si94, test_si95, test_si96, test_si97,
         test_si98, test_si99, test_si100;
  output g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435,
         g25442, g25489, g26104, g26135, g26149, g27380, g3993, g4088, g4090,
         g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549,
         g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738,
         g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518,
         g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944,
         g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334,
         g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012,
         g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249,
         g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266,
         g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275,
         test_so1, test_so2, test_so3, test_so4, test_so5, test_so6, test_so7,
         test_so8, test_so9, test_so10, test_so11, test_so12, test_so13,
         test_so14, test_so15, test_so16, test_so17, test_so18, test_so19,
         test_so20, test_so21, test_so22, test_so23, test_so24, test_so25,
         test_so26, test_so27, test_so28, test_so29, test_so30, test_so31,
         test_so32, test_so33, test_so34, test_so35, test_so36, test_so37,
         test_so38, test_so39, test_so40, test_so41, test_so42, test_so43,
         test_so44, test_so45, test_so46, test_so47, test_so48, test_so49,
         test_so50, test_so51, test_so52, test_so53, test_so54, test_so55,
         test_so56, test_so57, test_so58, test_so59, test_so60, test_so61,
         test_so62, test_so63, test_so64, test_so65, test_so66, test_so67,
         test_so68, test_so69, test_so70, test_so71, test_so72, test_so73,
         test_so74, test_so75, test_so76, test_so77, test_so78, test_so79,
         test_so80, test_so81, test_so82, test_so83, test_so84, test_so85,
         test_so86, test_so87, test_so88, test_so89, test_so90, test_so91,
         test_so92, test_so93, test_so94, test_so95, test_so96, test_so97,
         test_so98, test_so99, test_so100;
  wire   N690, N995, g2950, g2883, g2888, g2896, g2892, g2903, g2900, g2908,
         g2912, g2917, g2924, g2920, g2879, g2934, g2935, g2938, g2941, g2944,
         g2947, g2953, g2956, g2959, g2962, g2963, g2969, g2972, g2975, g2978,
         g2981, g2874, g1506, g1501, g1496, g1491, g1486, g1481, g1476, g1471,
         g2877, g8251, g813, g809, g805, g801, g797, g793, g789, g785, g7519,
         g2873, g125, g121, g117, g113, g109, g105, g101, g4450, g97, g2857,
         g2200, g2195, g2190, g2185, g2180, g2175, g2170, g2165, g2878, g3129,
         g3117, g3109, g3211, g3084, g3085, g3086, g3087, g3091, g3092, g3093,
         g3094, g3095, g3096, g3097, g3098, g3099, g3100, g3102, g3103, g3104,
         g3105, g3106, g3107, g3108, g3155, g3158, g3161, g3164, g3167, g3170,
         g3173, g3176, g3182, g3185, g3088, g3197, g3201, g3204, g3207, g3188,
         g3133, g3128, g3124, g3112, g3110, g3111, g3151, g3142, g185, g138,
         g165, g130, g131, g129, g133, g134, g132, g142, g143, g141, g145,
         g146, g148, g149, g147, g151, g152, g150, g154, g155, g153, g157,
         g158, g156, g160, g161, g159, g164, g162, g169, g170, g168, g172,
         g173, g171, g175, g176, g174, g178, g179, g177, g186, g192, g231,
         g234, g237, g195, g198, g201, g240, g243, g246, g204, g207, g210,
         g249, g252, g213, g216, g219, g258, g261, g264, g222, g225, g228,
         g267, g270, g273, g92, g88, g83, g74, g70, g65, g61, g56, g52, g180,
         g181, g276, g401, g309, g354, g343, g369, g358, g361, g384, g373,
         g376, g398, g388, g391, g408, g411, g414, g417, g420, g423, g428,
         g426, g429, g432, g435, g438, g441, g444, g448, g449, g447, g312,
         g313, g314, g315, g317, g318, g319, g320, g322, g323, g321, g403,
         g404, g402, g450, g452, g454, g280, g282, g284, g286, g288, g290,
         g305, g349, g350, g351, g352, g353, g357, g364, g365, g366, g367,
         g368, g372, g379, g380, g381, g383, g387, g394, g395, g396, g397,
         g324, g337, g545, g551, g550, g554, g557, g513, g523, g524, g564,
         g569, g570, g571, g572, g573, g574, g565, g566, g567, g568, g489,
         g7909, g485, g486, g487, g488, g455, g458, g461, g477, g478, g479,
         g480, g484, g464, g465, g471, g528, g535, g542, g543, g544, g548,
         g549, g499, g558, g559, g576, g577, g575, g579, g578, g582, g583,
         g581, g585, g586, g584, g587, g590, g593, g596, g599, g602, g614,
         g617, g605, g608, g611, g490, g493, g496, g506, g525, g536, g537,
         g538, g629, g630, g659, g640, g633, g653, g646, g660, g672, g679,
         g686, g692, g699, g700, g698, g702, g703, g701, g705, g706, g704,
         g708, g709, g707, g712, g710, g714, g715, g713, g717, g718, g716,
         g720, g721, g719, g723, g724, g722, g726, g725, g729, g730, g728,
         g732, g733, g731, g735, g736, g734, g738, g739, g737, g818, g819,
         g817, g821, g822, g820, g830, g831, g829, g833, g834, g832, g836,
         g837, g835, g840, g838, g842, g843, g841, g845, g846, g844, g848,
         g849, g847, g851, g852, g850, g857, g856, g860, g861, g859, g863,
         g864, g862, g866, g867, g865, g873, g876, g879, g918, g921, g882,
         g885, g888, g927, g930, g933, g891, g894, g897, g936, g939, g942,
         g900, g903, g906, g948, g951, g909, g912, g915, g954, g957, g960,
         g780, g776, g771, g767, g762, g758, g753, g744, g740, g868, g869,
         g963, g1092, g1088, g996, g1041, g1030, g1033, g1056, g1045, g1048,
         g1060, g1063, g1085, g1075, g1078, g1095, g1098, g1101, g1104, g1107,
         g1110, g1114, g1115, g1113, g1116, g1122, g1125, g1128, g1131, g1135,
         g1136, g1134, g999, g1000, g1001, g1002, g1003, g1004, g1005, g1006,
         g1009, g1010, g1008, g1090, g1091, g1089, g1137, g1139, g1141, g967,
         g969, g971, g973, g975, g977, g986, g992, g1029, g1036, g1037, g1038,
         g1040, g1044, g1051, g1052, g1053, g1054, g1055, g1059, g1066, g1067,
         g1068, g1069, g1070, g1074, g1081, g1083, g1084, g1011, g1024, g1231,
         g1237, g1236, g1240, g1243, g1196, g1199, g1209, g1210, g1255, g1256,
         g1257, g1258, g1259, g1260, g1251, g1252, g1253, g1254, g1176, g1172,
         g1173, g1175, g1142, g1145, g1148, g1164, g1165, g1166, g1167, g1171,
         g1151, g1152, g1155, g1158, g1214, g1221, g1229, g1235, g1186, g1244,
         g1245, g1262, g1263, g1261, g1265, g1266, g1264, g1268, g1269, g1271,
         g1272, g1270, g1273, g1276, g1279, g1282, g1285, g1288, g1300, g1303,
         g1306, g1291, g1294, g1297, g1180, g1183, g1192, g1211, g1222, g1223,
         g1224, g1315, g1316, g1345, g1326, g1319, g1339, g1332, g1346, g1358,
         g1352, g1365, g1372, g1378, g1386, g1384, g1388, g1389, g1387, g1391,
         g1392, g1390, g1394, g1395, g1393, g1397, g1398, g1396, g1400, g1399,
         g1403, g1404, g1402, g1406, g1407, g1405, g1409, g1410, g1408, g1412,
         g1413, g1411, g1415, g1416, g1418, g1419, g1417, g1421, g1422, g1420,
         g1424, g1425, g1423, g1520, g1547, g1512, g1513, g1511, g1516, g1514,
         g1524, g1525, g1523, g1527, g1528, g1526, g1530, g1531, g1529, g1533,
         g1534, g1532, g1536, g1535, g1539, g1540, g1538, g1542, g1543, g1541,
         g1545, g1546, g1544, g1551, g1552, g1550, g1554, g1555, g1557, g1558,
         g1556, g1560, g1561, g1559, g1567, g1570, g1573, g1612, g1615, g1618,
         g1576, g1579, g1582, g1624, g1627, g1585, g1588, g1591, g1630, g1633,
         g1636, g1594, g1597, g1600, g1639, g1642, g1645, g1603, g1609, g1648,
         g1651, g1654, g1466, g1462, g1457, g1453, g1448, g1444, g1439, g1435,
         g1430, g1426, g1562, g5612, g1563, g1657, g1786, g1782, g1690, g1735,
         g1724, g1727, g1750, g1739, g1742, g1765, g1754, g1757, g1779, g1772,
         g1789, g1792, g1795, g1798, g1801, g1804, g1808, g1809, g1807, g1810,
         g1813, g1816, g1819, g1822, g1829, g1830, g1828, g1693, g1694, g1695,
         g1696, g1697, g1698, g1699, g1700, g1701, g1703, g1704, g1702, g1785,
         g1783, g1831, g1833, g1835, g1661, g1663, g1665, g1667, g1669, g1671,
         g1680, g1686, g1723, g1730, g1731, g1732, g1733, g1734, g1738, g1745,
         g1747, g1748, g1749, g1753, g1760, g1761, g1762, g1763, g1764, g1768,
         g1775, g1776, g1777, g1778, g1705, g5695, g1718, g1925, g1931, g1930,
         g1934, g1937, g1890, g1893, g1903, g1904, g1944, g1949, g1950, g1951,
         g1953, g1954, g1945, g1946, g1947, g1948, g1870, g1866, g1867, g1868,
         g1869, g1836, g1842, g1858, g1859, g1860, g1861, g1865, g1845, g1846,
         g1849, g1852, g1908, g1915, g1922, g1923, g1929, g1880, g1938, g1939,
         g1956, g1957, g1955, g1959, g1960, g1958, g1962, g1963, g1961, g1966,
         g1964, g1967, g1970, g1973, g1976, g1979, g1982, g1994, g1997, g2000,
         g1985, g1988, g1991, g1874, g1877, g1886, g1905, g1916, g1917, g2009,
         g2010, g2039, g2020, g2013, g2033, g2026, g2040, g2052, g2046, g2059,
         g2072, g2079, g2080, g2078, g2082, g2083, g2081, g2085, g2086, g2084,
         g2088, g2089, g2087, g2091, g2090, g2094, g2095, g2093, g2097, g2098,
         g2096, g2100, g2101, g2099, g2103, g2104, g2102, g2106, g2105, g2109,
         g2110, g2108, g2112, g2113, g2111, g2115, g2116, g2114, g2118, g2119,
         g2117, g2214, g7084, g2241, g2206, g2207, g2205, g2209, g2210, g2208,
         g2218, g2219, g2217, g2221, g2222, g2220, g2224, g2223, g2227, g2228,
         g2226, g2230, g2231, g2229, g2233, g2234, g2232, g2236, g2237, g2235,
         g2239, g2238, g2245, g2246, g2244, g2248, g2249, g2247, g2251, g2252,
         g2250, g2254, g2255, g2253, g2261, g2267, g2306, g2309, g2312, g2270,
         g2273, g2276, g2315, g2318, g2321, g2279, g2282, g2285, g2324, g2330,
         g2288, g2291, g2294, g2333, g2336, g2339, g2297, g2300, g2303, g2342,
         g2345, g2348, g2160, g2151, g2147, g2142, g2138, g2133, g2129, g2124,
         g2120, g2256, g2257, g2351, g2480, g2476, g2429, g2418, g2421, g2444,
         g2433, g2436, g2459, g2448, g2451, g2473, g2463, g2466, g2483, g2486,
         g2492, g2495, g2498, g2502, g2503, g2501, g2504, g2507, g2510, g2513,
         g2516, g2519, g2523, g2524, g2387, g2388, g2389, g2390, g2391, g2392,
         g2393, g2394, g2395, g2397, g2398, g2396, g2478, g2479, g2525, g2527,
         g2529, g2355, g2357, g2359, g2361, g2365, g2374, g2380, g2417, g2424,
         g2425, g2426, g2427, g2428, g2432, g2439, g2441, g2442, g2443, g2447,
         g2454, g2455, g2456, g2457, g2458, g2462, g2469, g2470, g2471, g2472,
         g2412, g2619, g2625, g2624, g2628, g2631, g2584, g2587, g2597, g2598,
         g2638, g2643, g2645, g2646, g2647, g2648, g2639, g2640, g2641, g2642,
         g2564, g2560, g2561, g2562, g2530, g2533, g2536, g2552, g2553, g2554,
         g2555, g2559, g2539, g2540, g2543, g2546, g2602, g2609, g2617, g2623,
         g2574, g2632, g2633, g2650, g2651, g2649, g2653, g2654, g2652, g2656,
         g2655, g2659, g2660, g2658, g2661, g2664, g2667, g2670, g2673, g2676,
         g2688, g2691, g2694, g2679, g2685, g2565, g2568, g2571, g2580, g2599,
         g2611, g2612, g2703, g2704, g2733, g2714, g2707, g2727, g2720, g2734,
         g2746, g2753, g2760, g2766, g2773, g2774, g2772, g2776, g2777, g2775,
         g2779, g2780, g2778, g2782, g2783, g2785, g2786, g2784, g2788, g2789,
         g2787, g2791, g2792, g2790, g2794, g2795, g2793, g2797, g2798, g2800,
         g2801, g2799, g2803, g2804, g2802, g2806, g2807, g2805, g2809, g2810,
         g2808, g2812, g2813, g3080, g3043, g3044, g3045, g3046, g3047, g3048,
         g3049, g3050, g3051, g3052, g3053, g3056, g3057, g3058, g3059, g3060,
         g3061, g3062, g3063, g3064, g3065, g3066, g3067, g3068, g3069, g3071,
         g3072, g3073, g3074, g3075, g3076, g3077, g3078, g2997, g2993, g3006,
         g3002, g3013, g3024, g3018, g3028, g3036, g3032, g2987, g8270, g3083,
         g2990, g8258, g13149, g13111, g13155, g13160, g13124, g13164, g12487,
         g13171, g13135, g13175, g12507, g13182, g13143, g12524, g13194,
         g12457, g12539, g12467, g12482, g12499, g13110, g18669, g18678,
         g18707, g18719, g18726, g18743, g18755, g18763, g18780, g18782,
         g18794, g18821, g18804, g18820, g18835, g18852, g18836, g18975,
         g18837, g18866, g18968, g18883, g18867, g18868, g18885, g18754,
         g18906, g18907, g18781, g18803, g18942, g18957, g16654, g16671,
         g16692, g16718, g16860, g16866, g16803, g16824, g16835, g16844,
         g16845, g16851, g16853, g16854, g16857, g16861, g16880, g16802,
         g16823, g17222, g17224, g17225, g17226, g17228, g17229, g17234,
         g17235, g17236, g17246, g17247, g17248, g17269, g17270, g17271,
         g17302, g17303, g17340, g17341, g17383, g17429, g20310, g20314,
         g20333, g20343, g20353, g20375, g20376, g20417, g19144, g19149,
         g19153, g19154, g19157, g19162, g19163, g19167, g19172, g19173,
         g19178, g19184, g21842, g21843, g21845, g21847, g21851, g21878,
         g21880, g21882, g20874, g20875, g20876, g20879, g20880, g20881,
         g20882, g20883, g20682, g20891, g20892, g20893, g20894, g20896,
         g20897, g20898, g20899, g20900, g20901, g20902, g20903, g20717,
         g20910, g20911, g20912, g20913, g20915, g20916, g20917, g20918,
         g20919, g20921, g20922, g20923, g20924, g20925, g20926, g20927,
         g20752, g20934, g20935, g20936, g20937, g20939, g20940, g20941,
         g20944, g20945, g20946, g20947, g20948, g20949, g20950, g20951,
         g20952, g20953, g20954, g20955, g20789, g20962, g20963, g20964,
         g20965, g20966, g20967, g20968, g20969, g20970, g20972, g20973,
         g20974, g20975, g20976, g20977, g20978, g20979, g20980, g20981,
         g20982, g20983, g20989, g20990, g20991, g20992, g20993, g20994,
         g20995, g20996, g20997, g20999, g21000, g21001, g21002, g21003,
         g21004, g21005, g21006, g21007, g21009, g21010, g21011, g21015,
         g21016, g21017, g21018, g21019, g21020, g21021, g21022, g21023,
         g21025, g21026, g21027, g21028, g21029, g21031, g21032, g21033,
         g21034, g21035, g21039, g21040, g21041, g21042, g21043, g21044,
         g21045, g21046, g21047, g21051, g21052, g21053, g21054, g21055,
         g21056, g21060, g21061, g21062, g21063, g21070, g21071, g21072,
         g21073, g21074, g21075, g21080, g21081, g21082, g21094, g20877,
         g20884, g21346, g23000, g23117, g23014, g23126, g23022, g23030,
         g23137, g23039, g23047, g21970, g23058, g23067, g23076, g23081,
         g23092, g23093, g23097, g23110, g23111, g23114, g23123, g23124,
         g23132, g23133, g22025, g22027, g22028, g22029, g22030, g22031,
         g22032, g22033, g22034, g22035, g22037, g22038, g22039, g22040,
         g22041, g22042, g22043, g22044, g22045, g22047, g22048, g22049,
         g23136, g22054, g22055, g22056, g22057, g22058, g22059, g22060,
         g22061, g22063, g22064, g22065, g22066, g22067, g22068, g21969,
         g22073, g22074, g22075, g22076, g22077, g22078, g22079, g22080,
         g22081, g22087, g22088, g22089, g22090, g22091, g22092, g21972,
         g22097, g22098, g22099, g22100, g22101, g22102, g22103, g22104,
         g22105, g22106, g22112, g22113, g22114, g22115, g22116, g22117,
         g21974, g22122, g22123, g22124, g22125, g22126, g22127, g22128,
         g22129, g22130, g22131, g22132, g22138, g22139, g22140, g22141,
         g22142, g22143, g22145, g22146, g22147, g22148, g22149, g22150,
         g22151, g22152, g22153, g22154, g22155, g22161, g22162, g22163,
         g22164, g22166, g22167, g22168, g22169, g22170, g22171, g22172,
         g22173, g22177, g22178, g22179, g22180, g22182, g22183, g22184,
         g22185, g22191, g22192, g22193, g22194, g22200, g22578, g22615,
         g22651, g22026, g22218, g22687, g22231, g22234, g22242, g22247,
         g22249, g22263, g22267, g22269, g22280, g22284, g22299, g23399,
         g23406, g24174, g23413, g24178, g24179, g23418, g24181, g24182,
         g24206, g24207, g24208, g24209, g24212, g24213, g24214, g24215,
         g24216, g24218, g24219, g24222, g24223, g24225, g24226, g24228,
         g24230, g24231, g24235, g24237, g24238, g24243, g24250, g23385,
         g23392, g23400, g23324, g23407, g23329, g23330, g23339, g23348,
         g23357, g23358, g23359, g24059, g24072, g24083, g24092, g25027,
         g25042, g25056, g25067, g24426, g24430, g24434, g24438, g24491,
         g24498, g24499, g24501, g24507, g24508, g24510, g24511, g24513,
         g24445, g24446, g24519, g24521, g24522, g24524, g24525, g24527,
         g24532, g24534, g24535, g24537, g24538, g24545, g24547, g24548,
         g24557, g24473, g24476, g25932, g25935, g25938, g25940, g25204,
         g25206, g25207, g25209, g25211, g25212, g25213, g25214, g25215,
         g25217, g25218, g25219, g25220, g25221, g25222, g25223, g25224,
         g25225, g25227, g25228, g25229, g25230, g25231, g25232, g25233,
         g25234, g25235, g25236, g25237, g25239, g25240, g25241, g25242,
         g25243, g25244, g25245, g25246, g25247, g25248, g25249, g25250,
         g25251, g25252, g25253, g25185, g25255, g25256, g25257, g25189,
         g25259, g25265, g25191, g25260, g25194, g25262, g25263, g25197,
         g25266, g25267, g25268, g25270, g25271, g25272, g25279, g25280,
         g25199, g25288, g25201, g25202, g25450, g25451, g25452, g26541,
         g26545, g26547, g26553, g26557, g26559, g26569, g26573, g26575,
         g26592, g26596, g26616, g26529, g26530, g26655, g26531, g26659,
         g26661, g26532, g26664, g26665, g26667, g26669, g26670, g26672,
         g26675, g26676, g26025, g26660, g26666, g26671, g26677, g26048,
         g26031, g26037, g26183, g27120, g27123, g27129, g27131, g26803,
         g26804, g26805, g26806, g26807, g26808, g26776, g26809, g26810,
         g26811, g26812, g26813, g26814, g26781, g26815, g26816, g26817,
         g26786, g26818, g26820, g26821, g26789, g26822, g26823, g26824,
         g26825, g26826, g26795, g26827, g26798, g27594, g27603, g27612,
         g27621, g27672, g27678, g27682, g27243, g27253, g27255, g27256,
         g27257, g27258, g27259, g27260, g27261, g27262, g27263, g27264,
         g27265, g27266, g27267, g27268, g27269, g27270, g27271, g27272,
         g27273, g27274, g27275, g27276, g27277, g27278, g27279, g27280,
         g27281, g27282, g27283, g27284, g27285, g27286, g27287, g27288,
         g27289, g27290, g27291, g27292, g27293, g27294, g27295, g27296,
         g27297, g27298, g27299, g27300, g27301, g27302, g27303, g27304,
         g27305, g27306, g27307, g27308, g27309, g27310, g27311, g27312,
         g27313, g27314, g27315, g27316, g27317, g27318, g27319, g27320,
         g27321, g27322, g27323, g27324, g27325, g27326, g27327, g27328,
         g27329, g27330, g27331, g27332, g27333, g27334, g27335, g27336,
         g27337, g27338, g27339, g27340, g27341, g27342, g27343, g27344,
         g27345, g27346, g27347, g27348, g27354, g28145, g28146, g28147,
         g28148, g28199, g27718, g27722, g27724, g27759, g27760, g27761,
         g27762, g27763, g27764, g27765, g27766, g27767, g27768, g27769,
         g27771, g28634, g28635, g28636, g28637, g28668, g28321, g28325,
         g28328, g28342, g28344, g28345, g28346, g28348, g28349, g28350,
         g28351, g28352, g28353, g28354, g28355, g28356, g28357, g28358,
         g28360, g28361, g28362, g28363, g28364, g28366, g28367, g28368,
         g28371, g28420, g28421, g28425, g29109, g29110, g29111, g29112,
         g28732, g28735, g28736, g28738, g28744, g28745, g28746, g28747,
         g28749, g28754, g28758, g28759, g28760, g28761, g28990, g28763,
         g28767, g28771, g28772, g28773, g28774, g28778, g28782, g28783,
         g28788, g28903, g29353, g29354, g29355, g29357, g29167, g29169,
         g29170, g29172, g29173, g29178, g29179, g29181, g29182, g29184,
         g29185, g29187, g29194, g29197, g29198, g29201, g29204, g29205,
         g29209, g29212, g29213, g29218, g29221, g29226, g29579, g29606,
         g29608, g29580, g29609, g29611, g29612, g29581, g29613, g29616,
         g29617, g29582, g29618, g29620, g29621, g29623, g29936, g29939,
         g29941, g30055, g30072, g30061, g30267, g30268, g30269, g30270,
         g30271, g30272, g30273, g30274, g30275, g30276, g30277, g30278,
         g30279, g30280, g30281, g30282, g30283, g30284, g30285, g30286,
         g30287, g30288, g30289, g30290, g30291, g30292, g30293, g30294,
         g30295, g30296, g30297, g30298, g30299, g30300, g30301, g30302,
         g30303, g30304, g30245, g30246, g30247, g30248, g30249, g30250,
         g30251, g30252, g30253, g30254, g30255, g30256, g30257, g30258,
         g30259, g30260, g30261, g30262, g30263, g30264, g30265, g30266,
         g30455, g30468, g30470, g30482, g30485, g30487, g30500, g30503,
         g30505, g30338, g30341, g30356, g30668, g30669, g30670, g30671,
         g30672, g30673, g30674, g30675, g30676, g30677, g30678, g30679,
         g30680, g30681, g30682, g30683, g30684, g30686, g30687, g30688,
         g30689, g30690, g30691, g30692, g30693, g30694, g30695, g30699,
         g30700, g30701, g30702, g30703, g30704, g30705, g30706, g30707,
         g30708, g30709, g30566, g30635, g30636, g30637, g30638, g30639,
         g30640, g30641, g30642, g30643, g30644, g30645, g30646, g30647,
         g30648, g30649, g30650, g30651, g30652, g30653, g30654, g30655,
         g30656, g30657, g30658, g30659, g30660, g30661, g30662, g30663,
         g30664, g30665, g30666, g30667, g30796, g30798, g30801, DFF_1_n1,
         DFF_2_n1, DFF_15_n1, DFF_16_n1, DFF_18_n1, DFF_131_n1, DFF_132_n1,
         DFF_134_n1, DFF_140_n1, DFF_142_n1, DFF_144_n1, DFF_146_n1,
         DFF_149_n1, DFF_155_n1, DFF_156_n1, DFF_299_n1, DFF_301_n1,
         DFF_303_n1, DFF_305_n1, DFF_307_n1, DFF_309_n1, DFF_311_n1,
         DFF_313_n1, DFF_328_n1, DFF_444_n1, DFF_445_n1, DFF_446_n1,
         DFF_447_n1, DFF_448_n1, DFF_449_n1, DFF_453_n1, DFF_649_n1,
         DFF_651_n1, DFF_653_n1, DFF_655_n1, DFF_657_n1, DFF_659_n1,
         DFF_661_n1, DFF_663_n1, DFF_783_n1, DFF_792_n1, DFF_794_n1,
         DFF_795_n1, DFF_796_n1, DFF_797_n1, DFF_798_n1, DFF_799_n1,
         DFF_803_n1, DFF_999_n1, DFF_1001_n1, DFF_1003_n1, DFF_1005_n1,
         DFF_1007_n1, DFF_1009_n1, DFF_1011_n1, DFF_1013_n1, DFF_1099_n1,
         DFF_1100_n1, DFF_1133_n1, DFF_1142_n1, DFF_1144_n1, DFF_1145_n1,
         DFF_1146_n1, DFF_1147_n1, DFF_1148_n1, DFF_1149_n1, DFF_1153_n1,
         DFF_1349_n1, DFF_1351_n1, DFF_1353_n1, DFF_1355_n1, DFF_1357_n1,
         DFF_1359_n1, DFF_1361_n1, DFF_1363_n1, DFF_1378_n1, DFF_1449_n1,
         DFF_1450_n1, DFF_1494_n1, DFF_1495_n1, DFF_1496_n1, DFF_1497_n1,
         DFF_1498_n1, DFF_1499_n1, DFF_1503_n1, DFF_1561_n1, DFF_1562_n1,
         DFF_1612_n1, DFF_1616_n1, DFF_1617_n1, DFF_1618_n1, DFF_1625_n1,
         DFF_1626_n1, DFF_1628_n1, n1565, n1566, n1567, n1568, n1569, n1570,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1626, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1638, n1640, n1642, n1645, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1657, n1659, n1661, n1664,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1676, n1678, n1680,
         n1683, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1695, n1697,
         n1699, n1702, n1745, n1746, n1747, n1748, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1776, n1778, n1780, n1781, n1782, n1783, n1784, n1785, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1801, n1802, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1828, n1829, n1832, n1833, n1840, n1841, n1842,
         n1843, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1857, n1859, n1860, n1873, n1874, n1875, n1876, n1877,
         n1878, n1880, n1882, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1905, n1906, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1932, n1933, n1941, n1942, n1943, n1944, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1958,
         n1960, n1961, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1982,
         n1984, n1986, n1987, n1988, n1989, n1990, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2007,
         n2008, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2034, n2035,
         n2043, n2044, n2045, n2046, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2060, n2062, n2063, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2084, n2086, n2088, n2089, n2090,
         n2091, n2092, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2109, n2110, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2136, n2137, n2145, n2146, n2147, n2148,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2162, n2164, n2165, n2180, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3718, n3719, n3720, n3721, n3722, n3724, n3725, n3726, n3727, n3729,
         n3730, n3731, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3850, n3851, n3852, n3853, n3854, n3855, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4589, n4591, n4592, n4593, n4595,
         n4596, n4597, n4598, n4599, n4600, n4602, n4604, n4605, n4606, n4608,
         n4610, n4611, n4612, n4614, n4616, n4617, n4618, n4620, n4622, n4623,
         n4624, n4626, n4628, n4629, n4630, n4633, n4634, n4636, n4638, n4639,
         n4640, n4641, n4643, n4644, n4646, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n7907, n7909, n7912, n7913, n7918, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7929, n7930, n7936, n7937,
         n7938, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7960, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7971, n7978, n7979, n7980,
         n7983, n7984, n7985, n7986, n7987, n7988, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8017, n8018, n8019, n8020, n8021, n8024, n8025,
         n8026, n8027, n8040, n8043, n8044, n8045, n8046, n8047, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8065, n8066, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8086, n8087, n8088,
         n8089, n8090, n8098, n8099, n8102, n8103, n8104;
  assign test_so3 = g8251;
  assign test_so4 = g7519;
  assign test_so5 = g4450;
  assign test_so23 = g7909;
  assign test_so57 = g5612;
  assign test_so63 = g5695;
  assign test_so73 = g7084;
  assign test_so99 = g8270;
  assign test_so100 = g8258;

  LSDNENX1 U3772 ( .D(n2230), .ENB(n2217), .Q(n2231) );
  LSDNENX1 U3776 ( .D(n2374), .ENB(n2361), .Q(n2375) );
  LSDNENX1 U3777 ( .D(n4586), .ENB(DFF_2_n1), .Q(n4264) );
  LSDNENX1 U3778 ( .D(n2445), .ENB(n2446), .Q(n2440) );
  LSDNENX1 U3779 ( .D(n2478), .ENB(n2446), .Q(n2426) );
  LSDNENX1 U3780 ( .D(n2670), .ENB(n2671), .Q(n2669) );
  LSDNENX1 U3781 ( .D(n2685), .ENB(n2686), .Q(n2684) );
  LSDNENX1 U3782 ( .D(n2718), .ENB(n2719), .Q(n2717) );
  LSDNENX1 U3783 ( .D(n2982), .ENB(g2124), .Q(n2981) );
  LSDNENX1 U3784 ( .D(n2985), .ENB(g1430), .Q(n2984) );
  LSDNENX1 U3785 ( .D(n2988), .ENB(g744), .Q(n2987) );
  LSDNENX1 U3786 ( .D(n2991), .ENB(g56), .Q(n2990) );
  LSDNENX1 U3787 ( .D(n3742), .ENB(test_so98), .Q(n3741) );
  SDFFX1 DFF_0_Q_reg ( .D(n4586), .SI(test_si1), .SE(test_se), .CLK(CK), .Q(
        n8104), .QN(n1587) );
  SDFFX1 DFF_1_Q_reg ( .D(g16802), .SI(n8104), .SE(test_se), .CLK(CK), .Q(
        n8103), .QN(DFF_1_n1) );
  SDFFX1 DFF_2_Q_reg ( .D(g16823), .SI(n8103), .SE(test_se), .CLK(CK), .Q(
        n8102), .QN(DFF_2_n1) );
  SDFFX1 DFF_3_Q_reg ( .D(n4264), .SI(n8102), .SE(test_se), .CLK(CK), .Q(g2950), .QN(n4423) );
  SDFFX1 DFF_4_Q_reg ( .D(n4274), .SI(g2950), .SE(test_se), .CLK(CK), .Q(g2883), .QN(n4330) );
  SDFFX1 DFF_5_Q_reg ( .D(g22026), .SI(g2883), .SE(test_se), .CLK(CK), .Q(
        g2888), .QN() );
  SDFFX1 DFF_6_Q_reg ( .D(g23358), .SI(g2888), .SE(test_se), .CLK(CK), .Q(
        g2896), .QN(n4431) );
  SDFFX1 DFF_7_Q_reg ( .D(g24473), .SI(g2896), .SE(test_se), .CLK(CK), .Q(
        g2892), .QN() );
  SDFFX1 DFF_8_Q_reg ( .D(g25201), .SI(g2892), .SE(test_se), .CLK(CK), .Q(
        g2903), .QN(n4305) );
  SDFFX1 DFF_9_Q_reg ( .D(g26037), .SI(g2903), .SE(test_se), .CLK(CK), .Q(
        g2900), .QN(n4291) );
  SDFFX1 DFF_10_Q_reg ( .D(g26798), .SI(g2900), .SE(test_se), .CLK(CK), .Q(
        g2908), .QN(n4355) );
  SDFFX1 DFF_11_Q_reg ( .D(n4273), .SI(g2908), .SE(test_se), .CLK(CK), .Q(
        g2912), .QN(n4482) );
  SDFFX1 DFF_12_Q_reg ( .D(g23357), .SI(g2912), .SE(test_se), .CLK(CK), .Q(
        g2917), .QN(n4479) );
  SDFFX1 DFF_13_Q_reg ( .D(g24476), .SI(g2917), .SE(test_se), .CLK(CK), .Q(
        g2924), .QN(n4349) );
  SDFFX1 DFF_14_Q_reg ( .D(g25199), .SI(g2924), .SE(test_se), .CLK(CK), .Q(
        g2920), .QN() );
  SDFFX1 DFF_15_Q_reg ( .D(n4280), .SI(g2920), .SE(test_se), .CLK(CK), .Q(
        test_so1), .QN(DFF_15_n1) );
  SDFFX1 DFF_16_Q_reg ( .D(n4281), .SI(test_si2), .SE(test_se), .CLK(CK), .Q(
        n8099), .QN(DFF_16_n1) );
  SDFFX1 DFF_17_Q_reg ( .D(n4586), .SI(n8099), .SE(test_se), .CLK(CK), .Q(
        g8021), .QN() );
  SDFFX1 DFF_18_Q_reg ( .D(g8021), .SI(g8021), .SE(test_se), .CLK(CK), .Q(
        n8098), .QN(DFF_18_n1) );
  SDFFX1 DFF_19_Q_reg ( .D(n4279), .SI(n8098), .SE(test_se), .CLK(CK), .Q(
        g2879), .QN(n4351) );
  SDFFX1 DFF_20_Q_reg ( .D(g3212), .SI(g2879), .SE(test_se), .CLK(CK), .Q(
        g2934), .QN() );
  SDFFX1 DFF_21_Q_reg ( .D(g3228), .SI(g2934), .SE(test_se), .CLK(CK), .Q(
        g2935), .QN() );
  SDFFX1 DFF_22_Q_reg ( .D(g3227), .SI(g2935), .SE(test_se), .CLK(CK), .Q(
        g2938), .QN() );
  SDFFX1 DFF_23_Q_reg ( .D(g3226), .SI(g2938), .SE(test_se), .CLK(CK), .Q(
        g2941), .QN() );
  SDFFX1 DFF_24_Q_reg ( .D(g3225), .SI(g2941), .SE(test_se), .CLK(CK), .Q(
        g2944), .QN() );
  SDFFX1 DFF_25_Q_reg ( .D(g3224), .SI(g2944), .SE(test_se), .CLK(CK), .Q(
        g2947), .QN() );
  SDFFX1 DFF_26_Q_reg ( .D(g3223), .SI(g2947), .SE(test_se), .CLK(CK), .Q(
        g2953), .QN() );
  SDFFX1 DFF_27_Q_reg ( .D(g3222), .SI(g2953), .SE(test_se), .CLK(CK), .Q(
        g2956), .QN() );
  SDFFX1 DFF_28_Q_reg ( .D(g3221), .SI(g2956), .SE(test_se), .CLK(CK), .Q(
        g2959), .QN() );
  SDFFX1 DFF_29_Q_reg ( .D(g3232), .SI(g2959), .SE(test_se), .CLK(CK), .Q(
        g2962), .QN() );
  SDFFX1 DFF_30_Q_reg ( .D(g3220), .SI(g2962), .SE(test_se), .CLK(CK), .Q(
        g2963), .QN() );
  SDFFX1 DFF_31_Q_reg ( .D(g3219), .SI(g2963), .SE(test_se), .CLK(CK), .Q(
        test_so2), .QN() );
  SDFFX1 DFF_32_Q_reg ( .D(g3218), .SI(test_si3), .SE(test_se), .CLK(CK), .Q(
        g2969), .QN() );
  SDFFX1 DFF_33_Q_reg ( .D(g3217), .SI(g2969), .SE(test_se), .CLK(CK), .Q(
        g2972), .QN() );
  SDFFX1 DFF_34_Q_reg ( .D(g3216), .SI(g2972), .SE(test_se), .CLK(CK), .Q(
        g2975), .QN() );
  SDFFX1 DFF_35_Q_reg ( .D(g3215), .SI(g2975), .SE(test_se), .CLK(CK), .Q(
        g2978), .QN() );
  SDFFX1 DFF_36_Q_reg ( .D(g3214), .SI(g2978), .SE(test_se), .CLK(CK), .Q(
        g2981), .QN() );
  SDFFX1 DFF_37_Q_reg ( .D(g3213), .SI(g2981), .SE(test_se), .CLK(CK), .Q(
        g2874), .QN() );
  SDFFX1 DFF_38_Q_reg ( .D(g18754), .SI(g2874), .SE(test_se), .CLK(CK), .Q(
        g1506), .QN(n4288) );
  SDFFX1 DFF_39_Q_reg ( .D(g18781), .SI(g1506), .SE(test_se), .CLK(CK), .Q(
        g1501), .QN(n4565) );
  SDFFX1 DFF_40_Q_reg ( .D(g18803), .SI(g1501), .SE(test_se), .CLK(CK), .Q(
        g1496), .QN(n4557) );
  SDFFX1 DFF_41_Q_reg ( .D(g18821), .SI(g1496), .SE(test_se), .CLK(CK), .Q(
        g1491), .QN(n4326) );
  SDFFX1 DFF_42_Q_reg ( .D(g18835), .SI(g1491), .SE(test_se), .CLK(CK), .Q(
        g1486), .QN(n4390) );
  SDFFX1 DFF_43_Q_reg ( .D(g18852), .SI(g1486), .SE(test_se), .CLK(CK), .Q(
        g1481), .QN(n4320) );
  SDFFX1 DFF_44_Q_reg ( .D(g18866), .SI(g1481), .SE(test_se), .CLK(CK), .Q(
        g1476), .QN(n4374) );
  SDFFX1 DFF_45_Q_reg ( .D(g18883), .SI(g1476), .SE(test_se), .CLK(CK), .Q(
        g1471), .QN(n4378) );
  SDFFX1 DFF_46_Q_reg ( .D(g21880), .SI(g1471), .SE(test_se), .CLK(CK), .Q(
        g2877), .QN() );
  SDFFX1 DFF_47_Q_reg ( .D(g19154), .SI(g2877), .SE(test_se), .CLK(CK), .Q(
        g8251), .QN() );
  SDFFX1 DFF_48_Q_reg ( .D(g8251), .SI(test_si4), .SE(test_se), .CLK(CK), .Q(
        g813), .QN(n4289) );
  SDFFX1 DFF_49_Q_reg ( .D(g19163), .SI(g813), .SE(test_se), .CLK(CK), .Q(
        g4090), .QN() );
  SDFFX1 DFF_50_Q_reg ( .D(g4090), .SI(g4090), .SE(test_se), .CLK(CK), .Q(g809), .QN(n4567) );
  SDFFX1 DFF_51_Q_reg ( .D(g19173), .SI(g809), .SE(test_se), .CLK(CK), .Q(
        g4323), .QN() );
  SDFFX1 DFF_52_Q_reg ( .D(g4323), .SI(g4323), .SE(test_se), .CLK(CK), .Q(g805), .QN(n4559) );
  SDFFX1 DFF_53_Q_reg ( .D(g19184), .SI(g805), .SE(test_se), .CLK(CK), .Q(
        g4590), .QN() );
  SDFFX1 DFF_54_Q_reg ( .D(g4590), .SI(g4590), .SE(test_se), .CLK(CK), .Q(g801), .QN(n4327) );
  SDFFX1 DFF_55_Q_reg ( .D(g20310), .SI(g801), .SE(test_se), .CLK(CK), .Q(
        g6225), .QN() );
  SDFFX1 DFF_56_Q_reg ( .D(g6225), .SI(g6225), .SE(test_se), .CLK(CK), .Q(g797), .QN(n4391) );
  SDFFX1 DFF_57_Q_reg ( .D(g20343), .SI(g797), .SE(test_se), .CLK(CK), .Q(
        g6442), .QN() );
  SDFFX1 DFF_58_Q_reg ( .D(g6442), .SI(g6442), .SE(test_se), .CLK(CK), .Q(g793), .QN(n4321) );
  SDFFX1 DFF_59_Q_reg ( .D(g20376), .SI(g793), .SE(test_se), .CLK(CK), .Q(
        g6895), .QN() );
  SDFFX1 DFF_60_Q_reg ( .D(g6895), .SI(g6895), .SE(test_se), .CLK(CK), .Q(g789), .QN(n4375) );
  SDFFX1 DFF_61_Q_reg ( .D(g20417), .SI(g789), .SE(test_se), .CLK(CK), .Q(
        g7334), .QN() );
  SDFFX1 DFF_62_Q_reg ( .D(g7334), .SI(g7334), .SE(test_se), .CLK(CK), .Q(g785), .QN(n4379) );
  SDFFX1 DFF_63_Q_reg ( .D(g21878), .SI(g785), .SE(test_se), .CLK(CK), .Q(
        g7519), .QN() );
  SDFFX1 DFF_64_Q_reg ( .D(g7519), .SI(test_si5), .SE(test_se), .CLK(CK), .Q(
        g2873), .QN() );
  SDFFX1 DFF_65_Q_reg ( .D(g19153), .SI(g2873), .SE(test_se), .CLK(CK), .Q(
        g8249), .QN() );
  SDFFX1 DFF_66_Q_reg ( .D(g8249), .SI(g8249), .SE(test_se), .CLK(CK), .Q(g125), .QN(n4290) );
  SDFFX1 DFF_67_Q_reg ( .D(g19162), .SI(g125), .SE(test_se), .CLK(CK), .Q(
        g4088), .QN() );
  SDFFX1 DFF_68_Q_reg ( .D(g4088), .SI(g4088), .SE(test_se), .CLK(CK), .Q(g121), .QN(n4569) );
  SDFFX1 DFF_69_Q_reg ( .D(g19172), .SI(g121), .SE(test_se), .CLK(CK), .Q(
        g4321), .QN() );
  SDFFX1 DFF_70_Q_reg ( .D(g4321), .SI(g4321), .SE(test_se), .CLK(CK), .Q(g117), .QN(n4561) );
  SDFFX1 DFF_71_Q_reg ( .D(g19144), .SI(g117), .SE(test_se), .CLK(CK), .Q(
        g8023), .QN() );
  SDFFX1 DFF_72_Q_reg ( .D(g8023), .SI(g8023), .SE(test_se), .CLK(CK), .Q(g113), .QN(n4328) );
  SDFFX1 DFF_73_Q_reg ( .D(g19149), .SI(g113), .SE(test_se), .CLK(CK), .Q(
        g8175), .QN() );
  SDFFX1 DFF_74_Q_reg ( .D(g8175), .SI(g8175), .SE(test_se), .CLK(CK), .Q(g109), .QN(n4392) );
  SDFFX1 DFF_75_Q_reg ( .D(g19157), .SI(g109), .SE(test_se), .CLK(CK), .Q(
        g3993), .QN() );
  SDFFX1 DFF_76_Q_reg ( .D(g3993), .SI(g3993), .SE(test_se), .CLK(CK), .Q(g105), .QN(n4322) );
  SDFFX1 DFF_77_Q_reg ( .D(g19167), .SI(g105), .SE(test_se), .CLK(CK), .Q(
        g4200), .QN() );
  SDFFX1 DFF_78_Q_reg ( .D(g4200), .SI(g4200), .SE(test_se), .CLK(CK), .Q(g101), .QN(n4376) );
  SDFFX1 DFF_79_Q_reg ( .D(g19178), .SI(g101), .SE(test_se), .CLK(CK), .Q(
        g4450), .QN() );
  SDFFX1 DFF_80_Q_reg ( .D(g4450), .SI(test_si6), .SE(test_se), .CLK(CK), .Q(
        g97), .QN(n4380) );
  SDFFX1 DFF_81_Q_reg ( .D(g20874), .SI(g97), .SE(test_se), .CLK(CK), .Q(g8096), .QN() );
  SDFFX1 DFF_82_Q_reg ( .D(g8096), .SI(g8096), .SE(test_se), .CLK(CK), .Q(
        g2857), .QN() );
  SDFFX1 DFF_83_Q_reg ( .D(g18885), .SI(g2857), .SE(test_se), .CLK(CK), .Q(
        g2200), .QN(n4287) );
  SDFFX1 DFF_84_Q_reg ( .D(g18975), .SI(g2200), .SE(test_se), .CLK(CK), .Q(
        g2195), .QN(n4563) );
  SDFFX1 DFF_85_Q_reg ( .D(g18968), .SI(g2195), .SE(test_se), .CLK(CK), .Q(
        g2190), .QN(n4555) );
  SDFFX1 DFF_86_Q_reg ( .D(g18942), .SI(g2190), .SE(test_se), .CLK(CK), .Q(
        g2185), .QN(n4325) );
  SDFFX1 DFF_87_Q_reg ( .D(g18906), .SI(g2185), .SE(test_se), .CLK(CK), .Q(
        g2180), .QN(n4389) );
  SDFFX1 DFF_88_Q_reg ( .D(g18867), .SI(g2180), .SE(test_se), .CLK(CK), .Q(
        g2175), .QN(n4319) );
  SDFFX1 DFF_89_Q_reg ( .D(g18836), .SI(g2175), .SE(test_se), .CLK(CK), .Q(
        g2170), .QN(n4373) );
  SDFFX1 DFF_90_Q_reg ( .D(g18957), .SI(g2170), .SE(test_se), .CLK(CK), .Q(
        g2165), .QN(n4377) );
  SDFFX1 DFF_91_Q_reg ( .D(g21882), .SI(g2165), .SE(test_se), .CLK(CK), .Q(
        g2878), .QN() );
  SDFFX1 DFF_92_Q_reg ( .D(n4598), .SI(g2878), .SE(test_se), .CLK(CK), .Q(
        g3129), .QN(n4382) );
  SDFFX1 DFF_93_Q_reg ( .D(g8106), .SI(g3129), .SE(test_se), .CLK(CK), .Q(
        g3117), .QN(n4383) );
  SDFFX1 DFF_94_Q_reg ( .D(n4646), .SI(g3117), .SE(test_se), .CLK(CK), .Q(
        g3109), .QN(n4494) );
  SDFFX1 DFF_95_Q_reg ( .D(g18669), .SI(g3109), .SE(test_se), .CLK(CK), .Q(
        test_so6), .QN(n4446) );
  SDFFX1 DFF_96_Q_reg ( .D(g18719), .SI(test_si7), .SE(test_se), .CLK(CK), .Q(
        g3211), .QN(n4435) );
  SDFFX1 DFF_97_Q_reg ( .D(g18782), .SI(g3211), .SE(test_se), .CLK(CK), .Q(
        g3084), .QN(n4445) );
  SDFFX1 DFF_98_Q_reg ( .D(g17222), .SI(g3084), .SE(test_se), .CLK(CK), .Q(
        g3085), .QN(n4340) );
  SDFFX1 DFF_99_Q_reg ( .D(g17225), .SI(g3085), .SE(test_se), .CLK(CK), .Q(
        g3086), .QN(n4337) );
  SDFFX1 DFF_100_Q_reg ( .D(g17234), .SI(g3086), .SE(test_se), .CLK(CK), .Q(
        g3087), .QN(n4344) );
  SDFFX1 DFF_101_Q_reg ( .D(g17224), .SI(g3087), .SE(test_se), .CLK(CK), .Q(
        g3091), .QN(n4448) );
  SDFFX1 DFF_102_Q_reg ( .D(g17228), .SI(g3091), .SE(test_se), .CLK(CK), .Q(
        g3092), .QN(n4451) );
  SDFFX1 DFF_103_Q_reg ( .D(g17246), .SI(g3092), .SE(test_se), .CLK(CK), .Q(
        g3093), .QN(n4346) );
  SDFFX1 DFF_104_Q_reg ( .D(g17226), .SI(g3093), .SE(test_se), .CLK(CK), .Q(
        g3094), .QN(n4440) );
  SDFFX1 DFF_105_Q_reg ( .D(g17235), .SI(g3094), .SE(test_se), .CLK(CK), .Q(
        g3095), .QN(n4439) );
  SDFFX1 DFF_106_Q_reg ( .D(g17269), .SI(g3095), .SE(test_se), .CLK(CK), .Q(
        g3096), .QN(n4336) );
  SDFFX1 DFF_107_Q_reg ( .D(g25450), .SI(g3096), .SE(test_se), .CLK(CK), .Q(
        g3097), .QN(n4433) );
  SDFFX1 DFF_108_Q_reg ( .D(g25451), .SI(g3097), .SE(test_se), .CLK(CK), .Q(
        g3098), .QN(n4434) );
  SDFFX1 DFF_109_Q_reg ( .D(g25452), .SI(g3098), .SE(test_se), .CLK(CK), .Q(
        g3099), .QN(n4443) );
  SDFFX1 DFF_110_Q_reg ( .D(g28420), .SI(g3099), .SE(test_se), .CLK(CK), .Q(
        g3100), .QN(n4342) );
  SDFFX1 DFF_111_Q_reg ( .D(g28421), .SI(g3100), .SE(test_se), .CLK(CK), .Q(
        test_so7), .QN(n4335) );
  SDFFX1 DFF_112_Q_reg ( .D(g28425), .SI(test_si8), .SE(test_se), .CLK(CK), 
        .Q(g3102), .QN(n4343) );
  SDFFX1 DFF_113_Q_reg ( .D(g29936), .SI(g3102), .SE(test_se), .CLK(CK), .Q(
        g3103), .QN(n4447) );
  SDFFX1 DFF_114_Q_reg ( .D(g29939), .SI(g3103), .SE(test_se), .CLK(CK), .Q(
        g3104), .QN(n4452) );
  SDFFX1 DFF_115_Q_reg ( .D(g29941), .SI(g3104), .SE(test_se), .CLK(CK), .Q(
        g3105), .QN(n4347) );
  SDFFX1 DFF_116_Q_reg ( .D(g30796), .SI(g3105), .SE(test_se), .CLK(CK), .Q(
        g3106), .QN(n4438) );
  SDFFX1 DFF_117_Q_reg ( .D(g30798), .SI(g3106), .SE(test_se), .CLK(CK), .Q(
        g3107), .QN(n4437) );
  SDFFX1 DFF_118_Q_reg ( .D(g30801), .SI(g3107), .SE(test_se), .CLK(CK), .Q(
        g3108), .QN(n4334) );
  SDFFX1 DFF_119_Q_reg ( .D(g17229), .SI(g3108), .SE(test_se), .CLK(CK), .Q(
        g3155), .QN(n4449) );
  SDFFX1 DFF_120_Q_reg ( .D(g17247), .SI(g3155), .SE(test_se), .CLK(CK), .Q(
        g3158), .QN(n4436) );
  SDFFX1 DFF_121_Q_reg ( .D(g17302), .SI(g3158), .SE(test_se), .CLK(CK), .Q(
        g3161), .QN(n4444) );
  SDFFX1 DFF_122_Q_reg ( .D(g17236), .SI(g3161), .SE(test_se), .CLK(CK), .Q(
        g3164), .QN(n4339) );
  SDFFX1 DFF_123_Q_reg ( .D(g17270), .SI(g3164), .SE(test_se), .CLK(CK), .Q(
        g3167), .QN(n4348) );
  SDFFX1 DFF_124_Q_reg ( .D(g17340), .SI(g3167), .SE(test_se), .CLK(CK), .Q(
        g3170), .QN(n4441) );
  SDFFX1 DFF_125_Q_reg ( .D(g17248), .SI(g3170), .SE(test_se), .CLK(CK), .Q(
        g3173), .QN(n4338) );
  SDFFX1 DFF_126_Q_reg ( .D(g17303), .SI(g3173), .SE(test_se), .CLK(CK), .Q(
        g3176), .QN(n4450) );
  SDFFX1 DFF_127_Q_reg ( .D(g17383), .SI(g3176), .SE(test_se), .CLK(CK), .Q(
        test_so8), .QN(n4345) );
  SDFFX1 DFF_128_Q_reg ( .D(g17271), .SI(test_si9), .SE(test_se), .CLK(CK), 
        .Q(g3182), .QN(n4453) );
  SDFFX1 DFF_129_Q_reg ( .D(g17341), .SI(g3182), .SE(test_se), .CLK(CK), .Q(
        g3185), .QN(n4442) );
  SDFFX1 DFF_130_Q_reg ( .D(g17429), .SI(g3185), .SE(test_se), .CLK(CK), .Q(
        g3088), .QN(n4341) );
  SDFFX1 DFF_131_Q_reg ( .D(g24734), .SI(g3088), .SE(test_se), .CLK(CK), .Q(
        n8090), .QN(DFF_131_n1) );
  SDFFX1 DFF_132_Q_reg ( .D(g25442), .SI(n8090), .SE(test_se), .CLK(CK), .Q(
        n8089), .QN(DFF_132_n1) );
  SDFFX1 DFF_133_Q_reg ( .D(g25435), .SI(n8089), .SE(test_se), .CLK(CK), .Q(
        g3197), .QN() );
  SDFFX1 DFF_134_Q_reg ( .D(g25420), .SI(g3197), .SE(test_se), .CLK(CK), .Q(
        n8088), .QN(DFF_134_n1) );
  SDFFX1 DFF_135_Q_reg ( .D(g26149), .SI(n8088), .SE(test_se), .CLK(CK), .Q(
        g3201), .QN(n4406) );
  SDFFX1 DFF_136_Q_reg ( .D(g26135), .SI(g3201), .SE(test_se), .CLK(CK), .Q(
        g3204), .QN() );
  SDFFX1 DFF_137_Q_reg ( .D(g26104), .SI(g3204), .SE(test_se), .CLK(CK), .Q(
        g3207), .QN(n4329) );
  SDFFX1 DFF_138_Q_reg ( .D(g27380), .SI(g3207), .SE(test_se), .CLK(CK), .Q(
        g3188), .QN(n4405) );
  SDFFX1 DFF_139_Q_reg ( .D(n1576), .SI(g3188), .SE(test_se), .CLK(CK), .Q(
        g3133), .QN() );
  SDFFX1 DFF_140_Q_reg ( .D(g26104), .SI(g3133), .SE(test_se), .CLK(CK), .Q(
        n8087), .QN(DFF_140_n1) );
  SDFFX1 DFF_141_Q_reg ( .D(n1575), .SI(n8087), .SE(test_se), .CLK(CK), .Q(
        g3128), .QN() );
  SDFFX1 DFF_142_Q_reg ( .D(g26149), .SI(g3128), .SE(test_se), .CLK(CK), .Q(
        n8086), .QN(DFF_142_n1) );
  SDFFX1 DFF_143_Q_reg ( .D(g25420), .SI(n8086), .SE(test_se), .CLK(CK), .Q(
        test_so9), .QN() );
  SDFFX1 DFF_144_Q_reg ( .D(n1573), .SI(test_si10), .SE(test_se), .CLK(CK), 
        .Q(n8084), .QN(DFF_144_n1) );
  SDFFX1 DFF_145_Q_reg ( .D(g25442), .SI(n8084), .SE(test_se), .CLK(CK), .Q(
        g3124), .QN() );
  SDFFX1 DFF_146_Q_reg ( .D(n1572), .SI(g3124), .SE(test_se), .CLK(CK), .Q(
        n8083), .QN(DFF_146_n1) );
  SDFFX1 DFF_147_Q_reg ( .D(g26104), .SI(n8083), .SE(test_se), .CLK(CK), .Q(
        n8082), .QN(n4302) );
  SDFFX1 DFF_148_Q_reg ( .D(g26135), .SI(n8082), .SE(test_se), .CLK(CK), .Q(
        n8081), .QN(n4331) );
  SDFFX1 DFF_149_Q_reg ( .D(g26149), .SI(n8081), .SE(test_se), .CLK(CK), .Q(
        n8080), .QN(DFF_149_n1) );
  SDFFX1 DFF_150_Q_reg ( .D(g25420), .SI(n8080), .SE(test_se), .CLK(CK), .Q(
        g3112), .QN() );
  SDFFX1 DFF_151_Q_reg ( .D(g25435), .SI(g3112), .SE(test_se), .CLK(CK), .Q(
        g3110), .QN() );
  SDFFX1 DFF_152_Q_reg ( .D(g25442), .SI(g3110), .SE(test_se), .CLK(CK), .Q(
        g3111), .QN() );
  SDFFX1 DFF_153_Q_reg ( .D(g27380), .SI(g3111), .SE(test_se), .CLK(CK), .Q(
        n8079), .QN(n4425) );
  SDFFX1 DFF_154_Q_reg ( .D(g26104), .SI(n8079), .SE(test_se), .CLK(CK), .Q(
        n8078), .QN(n4332) );
  SDFFX1 DFF_155_Q_reg ( .D(g26135), .SI(n8078), .SE(test_se), .CLK(CK), .Q(
        n8077), .QN(DFF_155_n1) );
  SDFFX1 DFF_156_Q_reg ( .D(g26149), .SI(n8077), .SE(test_se), .CLK(CK), .Q(
        n8076), .QN(DFF_156_n1) );
  SDFFX1 DFF_157_Q_reg ( .D(g27380), .SI(n8076), .SE(test_se), .CLK(CK), .Q(
        g3151), .QN(n4424) );
  SDFFX1 DFF_158_Q_reg ( .D(g26104), .SI(g3151), .SE(test_se), .CLK(CK), .Q(
        g3142), .QN(n4301) );
  SDFFX1 DFF_159_Q_reg ( .D(g26135), .SI(g3142), .SE(test_se), .CLK(CK), .Q(
        test_so10), .QN(n4333) );
  SDFFX1 DFF_160_Q_reg ( .D(n1576), .SI(test_si11), .SE(test_se), .CLK(CK), 
        .Q(g185), .QN(n4384) );
  SDFFX1 DFF_161_Q_reg ( .D(n4650), .SI(g185), .SE(test_se), .CLK(CK), .Q(g138), .QN(n4318) );
  SDFFX1 DFF_162_Q_reg ( .D(g6231), .SI(g138), .SE(test_se), .CLK(CK), .Q(
        g6313), .QN(n4512) );
  SDFFX1 DFF_163_Q_reg ( .D(n4593), .SI(g6313), .SE(test_se), .CLK(CK), .Q(
        g165), .QN(n4369) );
  SDFFX1 DFF_164_Q_reg ( .D(g22100), .SI(g165), .SE(test_se), .CLK(CK), .Q(
        g130), .QN() );
  SDFFX1 DFF_165_Q_reg ( .D(g22122), .SI(g130), .SE(test_se), .CLK(CK), .Q(
        g131), .QN() );
  SDFFX1 DFF_166_Q_reg ( .D(g22141), .SI(g131), .SE(test_se), .CLK(CK), .Q(
        g129), .QN() );
  SDFFX1 DFF_167_Q_reg ( .D(g22123), .SI(g129), .SE(test_se), .CLK(CK), .Q(
        g133), .QN() );
  SDFFX1 DFF_168_Q_reg ( .D(g22142), .SI(g133), .SE(test_se), .CLK(CK), .Q(
        g134), .QN() );
  SDFFX1 DFF_169_Q_reg ( .D(g22161), .SI(g134), .SE(test_se), .CLK(CK), .Q(
        g132), .QN() );
  SDFFX1 DFF_170_Q_reg ( .D(g22025), .SI(g132), .SE(test_se), .CLK(CK), .Q(
        g142), .QN() );
  SDFFX1 DFF_171_Q_reg ( .D(g22027), .SI(g142), .SE(test_se), .CLK(CK), .Q(
        g143), .QN() );
  SDFFX1 DFF_172_Q_reg ( .D(g22030), .SI(g143), .SE(test_se), .CLK(CK), .Q(
        g141), .QN() );
  SDFFX1 DFF_173_Q_reg ( .D(g22028), .SI(g141), .SE(test_se), .CLK(CK), .Q(
        g145), .QN() );
  SDFFX1 DFF_174_Q_reg ( .D(g22031), .SI(g145), .SE(test_se), .CLK(CK), .Q(
        g146), .QN() );
  SDFFX1 DFF_175_Q_reg ( .D(g22037), .SI(g146), .SE(test_se), .CLK(CK), .Q(
        test_so11), .QN() );
  SDFFX1 DFF_176_Q_reg ( .D(g22032), .SI(test_si12), .SE(test_se), .CLK(CK), 
        .Q(g148), .QN() );
  SDFFX1 DFF_177_Q_reg ( .D(g22038), .SI(g148), .SE(test_se), .CLK(CK), .Q(
        g149), .QN() );
  SDFFX1 DFF_178_Q_reg ( .D(g22047), .SI(g149), .SE(test_se), .CLK(CK), .Q(
        g147), .QN() );
  SDFFX1 DFF_179_Q_reg ( .D(g22039), .SI(g147), .SE(test_se), .CLK(CK), .Q(
        g151), .QN() );
  SDFFX1 DFF_180_Q_reg ( .D(g22048), .SI(g151), .SE(test_se), .CLK(CK), .Q(
        g152), .QN() );
  SDFFX1 DFF_181_Q_reg ( .D(g22063), .SI(g152), .SE(test_se), .CLK(CK), .Q(
        g150), .QN() );
  SDFFX1 DFF_182_Q_reg ( .D(g22049), .SI(g150), .SE(test_se), .CLK(CK), .Q(
        g154), .QN() );
  SDFFX1 DFF_183_Q_reg ( .D(g22064), .SI(g154), .SE(test_se), .CLK(CK), .Q(
        g155), .QN() );
  SDFFX1 DFF_184_Q_reg ( .D(g22079), .SI(g155), .SE(test_se), .CLK(CK), .Q(
        g153), .QN() );
  SDFFX1 DFF_185_Q_reg ( .D(g22065), .SI(g153), .SE(test_se), .CLK(CK), .Q(
        g157), .QN() );
  SDFFX1 DFF_186_Q_reg ( .D(g22080), .SI(g157), .SE(test_se), .CLK(CK), .Q(
        g158), .QN() );
  SDFFX1 DFF_187_Q_reg ( .D(g22101), .SI(g158), .SE(test_se), .CLK(CK), .Q(
        g156), .QN() );
  SDFFX1 DFF_188_Q_reg ( .D(g22081), .SI(g156), .SE(test_se), .CLK(CK), .Q(
        g160), .QN() );
  SDFFX1 DFF_189_Q_reg ( .D(g22102), .SI(g160), .SE(test_se), .CLK(CK), .Q(
        g161), .QN() );
  SDFFX1 DFF_190_Q_reg ( .D(g22124), .SI(g161), .SE(test_se), .CLK(CK), .Q(
        g159), .QN() );
  SDFFX1 DFF_191_Q_reg ( .D(g22103), .SI(g159), .SE(test_se), .CLK(CK), .Q(
        test_so12), .QN() );
  SDFFX1 DFF_192_Q_reg ( .D(g22125), .SI(test_si13), .SE(test_se), .CLK(CK), 
        .Q(g164), .QN() );
  SDFFX1 DFF_193_Q_reg ( .D(g22143), .SI(g164), .SE(test_se), .CLK(CK), .Q(
        g162), .QN() );
  SDFFX1 DFF_194_Q_reg ( .D(g25204), .SI(g162), .SE(test_se), .CLK(CK), .Q(
        g169), .QN() );
  SDFFX1 DFF_195_Q_reg ( .D(g25206), .SI(g169), .SE(test_se), .CLK(CK), .Q(
        g170), .QN() );
  SDFFX1 DFF_196_Q_reg ( .D(g25211), .SI(g170), .SE(test_se), .CLK(CK), .Q(
        g168), .QN() );
  SDFFX1 DFF_197_Q_reg ( .D(g25207), .SI(g168), .SE(test_se), .CLK(CK), .Q(
        g172), .QN() );
  SDFFX1 DFF_198_Q_reg ( .D(g25212), .SI(g172), .SE(test_se), .CLK(CK), .Q(
        g173), .QN() );
  SDFFX1 DFF_199_Q_reg ( .D(g25218), .SI(g173), .SE(test_se), .CLK(CK), .Q(
        g171), .QN() );
  SDFFX1 DFF_200_Q_reg ( .D(g25213), .SI(g171), .SE(test_se), .CLK(CK), .Q(
        g175), .QN() );
  SDFFX1 DFF_201_Q_reg ( .D(g25219), .SI(g175), .SE(test_se), .CLK(CK), .Q(
        g176), .QN() );
  SDFFX1 DFF_202_Q_reg ( .D(g25228), .SI(g176), .SE(test_se), .CLK(CK), .Q(
        g174), .QN() );
  SDFFX1 DFF_203_Q_reg ( .D(g25220), .SI(g174), .SE(test_se), .CLK(CK), .Q(
        g178), .QN() );
  SDFFX1 DFF_204_Q_reg ( .D(g25229), .SI(g178), .SE(test_se), .CLK(CK), .Q(
        g179), .QN() );
  SDFFX1 DFF_205_Q_reg ( .D(g25239), .SI(g179), .SE(test_se), .CLK(CK), .Q(
        g177), .QN() );
  SDFFX1 DFF_206_Q_reg ( .D(g30261), .SI(g177), .SE(test_se), .CLK(CK), .Q(
        g186), .QN() );
  SDFFX1 DFF_207_Q_reg ( .D(g30267), .SI(g186), .SE(test_se), .CLK(CK), .Q(
        test_so13), .QN() );
  SDFFX1 DFF_208_Q_reg ( .D(g30275), .SI(test_si14), .SE(test_se), .CLK(CK), 
        .Q(g192), .QN() );
  SDFFX1 DFF_209_Q_reg ( .D(g30637), .SI(g192), .SE(test_se), .CLK(CK), .Q(
        g231), .QN() );
  SDFFX1 DFF_210_Q_reg ( .D(g30640), .SI(g231), .SE(test_se), .CLK(CK), .Q(
        g234), .QN() );
  SDFFX1 DFF_211_Q_reg ( .D(g30645), .SI(g234), .SE(test_se), .CLK(CK), .Q(
        g237), .QN() );
  SDFFX1 DFF_212_Q_reg ( .D(g30668), .SI(g237), .SE(test_se), .CLK(CK), .Q(
        g195), .QN() );
  SDFFX1 DFF_213_Q_reg ( .D(g30674), .SI(g195), .SE(test_se), .CLK(CK), .Q(
        g198), .QN() );
  SDFFX1 DFF_214_Q_reg ( .D(g30680), .SI(g198), .SE(test_se), .CLK(CK), .Q(
        g201), .QN() );
  SDFFX1 DFF_215_Q_reg ( .D(g30641), .SI(g201), .SE(test_se), .CLK(CK), .Q(
        g240), .QN() );
  SDFFX1 DFF_216_Q_reg ( .D(g30646), .SI(g240), .SE(test_se), .CLK(CK), .Q(
        g243), .QN() );
  SDFFX1 DFF_217_Q_reg ( .D(g30653), .SI(g243), .SE(test_se), .CLK(CK), .Q(
        g246), .QN() );
  SDFFX1 DFF_218_Q_reg ( .D(g30276), .SI(g246), .SE(test_se), .CLK(CK), .Q(
        g204), .QN() );
  SDFFX1 DFF_219_Q_reg ( .D(g30284), .SI(g204), .SE(test_se), .CLK(CK), .Q(
        g207), .QN() );
  SDFFX1 DFF_220_Q_reg ( .D(g30292), .SI(g207), .SE(test_se), .CLK(CK), .Q(
        g210), .QN() );
  SDFFX1 DFF_221_Q_reg ( .D(g30254), .SI(g210), .SE(test_se), .CLK(CK), .Q(
        g249), .QN() );
  SDFFX1 DFF_222_Q_reg ( .D(g30257), .SI(g249), .SE(test_se), .CLK(CK), .Q(
        g252), .QN() );
  SDFFX1 DFF_223_Q_reg ( .D(g30262), .SI(g252), .SE(test_se), .CLK(CK), .Q(
        test_so14), .QN() );
  SDFFX1 DFF_224_Q_reg ( .D(g30245), .SI(test_si15), .SE(test_se), .CLK(CK), 
        .Q(g213), .QN() );
  SDFFX1 DFF_225_Q_reg ( .D(g30246), .SI(g213), .SE(test_se), .CLK(CK), .Q(
        g216), .QN() );
  SDFFX1 DFF_226_Q_reg ( .D(g30248), .SI(g216), .SE(test_se), .CLK(CK), .Q(
        g219), .QN() );
  SDFFX1 DFF_227_Q_reg ( .D(g30258), .SI(g219), .SE(test_se), .CLK(CK), .Q(
        g258), .QN() );
  SDFFX1 DFF_228_Q_reg ( .D(g30263), .SI(g258), .SE(test_se), .CLK(CK), .Q(
        g261), .QN() );
  SDFFX1 DFF_229_Q_reg ( .D(g30268), .SI(g261), .SE(test_se), .CLK(CK), .Q(
        g264), .QN() );
  SDFFX1 DFF_230_Q_reg ( .D(g30635), .SI(g264), .SE(test_se), .CLK(CK), .Q(
        g222), .QN() );
  SDFFX1 DFF_231_Q_reg ( .D(g30636), .SI(g222), .SE(test_se), .CLK(CK), .Q(
        g225), .QN() );
  SDFFX1 DFF_232_Q_reg ( .D(g30639), .SI(g225), .SE(test_se), .CLK(CK), .Q(
        g228), .QN() );
  SDFFX1 DFF_233_Q_reg ( .D(g30661), .SI(g228), .SE(test_se), .CLK(CK), .Q(
        g267), .QN() );
  SDFFX1 DFF_234_Q_reg ( .D(g30669), .SI(g267), .SE(test_se), .CLK(CK), .Q(
        g270), .QN() );
  SDFFX1 DFF_235_Q_reg ( .D(g30675), .SI(g270), .SE(test_se), .CLK(CK), .Q(
        g273), .QN() );
  SDFFX1 DFF_236_Q_reg ( .D(g25027), .SI(g273), .SE(test_se), .CLK(CK), .Q(g92), .QN() );
  SDFFX1 DFF_237_Q_reg ( .D(g25932), .SI(g92), .SE(test_se), .CLK(CK), .Q(g88), 
        .QN() );
  SDFFX1 DFF_238_Q_reg ( .D(g26529), .SI(g88), .SE(test_se), .CLK(CK), .Q(g83), 
        .QN() );
  SDFFX1 DFF_239_Q_reg ( .D(g27120), .SI(g83), .SE(test_se), .CLK(CK), .Q(
        test_so15), .QN() );
  SDFFX1 DFF_240_Q_reg ( .D(g27594), .SI(test_si16), .SE(test_se), .CLK(CK), 
        .Q(g74), .QN() );
  SDFFX1 DFF_241_Q_reg ( .D(g28145), .SI(g74), .SE(test_se), .CLK(CK), .Q(g70), 
        .QN() );
  SDFFX1 DFF_242_Q_reg ( .D(g28634), .SI(g70), .SE(test_se), .CLK(CK), .Q(g65), 
        .QN() );
  SDFFX1 DFF_243_Q_reg ( .D(g29109), .SI(g65), .SE(test_se), .CLK(CK), .Q(g61), 
        .QN() );
  SDFFX1 DFF_244_Q_reg ( .D(g29353), .SI(g61), .SE(test_se), .CLK(CK), .Q(g56), 
        .QN() );
  SDFFX1 DFF_245_Q_reg ( .D(g29579), .SI(g56), .SE(test_se), .CLK(CK), .Q(g52), 
        .QN() );
  SDFFX1 DFF_246_Q_reg ( .D(g13110), .SI(g52), .SE(test_se), .CLK(CK), .Q(g180), .QN() );
  SDFFX1 DFF_247_Q_reg ( .D(g180), .SI(g180), .SE(test_se), .CLK(CK), .Q(g5549), .QN() );
  SDFFX1 DFF_248_Q_reg ( .D(g5549), .SI(g5549), .SE(test_se), .CLK(CK), .Q(
        g181), .QN() );
  SDFFX1 DFF_251_Q_reg ( .D(n4641), .SI(g6447), .SE(test_se), .CLK(CK), .Q(
        g401), .QN(n4506) );
  SDFFX1 DFF_252_Q_reg ( .D(g5549), .SI(g401), .SE(test_se), .CLK(CK), .Q(g309), .QN(n4388) );
  SDFFX1 DFF_253_Q_reg ( .D(g27253), .SI(g309), .SE(test_se), .CLK(CK), .Q(
        g354), .QN() );
  SDFFX1 DFF_254_Q_reg ( .D(g27255), .SI(g354), .SE(test_se), .CLK(CK), .Q(
        g343), .QN() );
  SDFFX1 DFF_255_Q_reg ( .D(g27258), .SI(g343), .SE(test_se), .CLK(CK), .Q(
        test_so16), .QN() );
  SDFFX1 DFF_256_Q_reg ( .D(g27256), .SI(test_si17), .SE(test_se), .CLK(CK), 
        .Q(g369), .QN() );
  SDFFX1 DFF_257_Q_reg ( .D(g27259), .SI(g369), .SE(test_se), .CLK(CK), .Q(
        g358), .QN() );
  SDFFX1 DFF_258_Q_reg ( .D(g27265), .SI(g358), .SE(test_se), .CLK(CK), .Q(
        g361), .QN() );
  SDFFX1 DFF_259_Q_reg ( .D(g27260), .SI(g361), .SE(test_se), .CLK(CK), .Q(
        g384), .QN() );
  SDFFX1 DFF_260_Q_reg ( .D(g27266), .SI(g384), .SE(test_se), .CLK(CK), .Q(
        g373), .QN() );
  SDFFX1 DFF_261_Q_reg ( .D(g27277), .SI(g373), .SE(test_se), .CLK(CK), .Q(
        g376), .QN() );
  SDFFX1 DFF_262_Q_reg ( .D(g27267), .SI(g376), .SE(test_se), .CLK(CK), .Q(
        g398), .QN() );
  SDFFX1 DFF_263_Q_reg ( .D(g27278), .SI(g398), .SE(test_se), .CLK(CK), .Q(
        g388), .QN() );
  SDFFX1 DFF_264_Q_reg ( .D(g27293), .SI(g388), .SE(test_se), .CLK(CK), .Q(
        g391), .QN() );
  SDFFX1 DFF_265_Q_reg ( .D(g28732), .SI(g391), .SE(test_se), .CLK(CK), .Q(
        g408), .QN() );
  SDFFX1 DFF_266_Q_reg ( .D(g28735), .SI(g408), .SE(test_se), .CLK(CK), .Q(
        g411), .QN() );
  SDFFX1 DFF_267_Q_reg ( .D(g28744), .SI(g411), .SE(test_se), .CLK(CK), .Q(
        g414), .QN() );
  SDFFX1 DFF_268_Q_reg ( .D(g29194), .SI(g414), .SE(test_se), .CLK(CK), .Q(
        g417), .QN() );
  SDFFX1 DFF_269_Q_reg ( .D(g29197), .SI(g417), .SE(test_se), .CLK(CK), .Q(
        g420), .QN() );
  SDFFX1 DFF_270_Q_reg ( .D(g29201), .SI(g420), .SE(test_se), .CLK(CK), .Q(
        g423), .QN() );
  SDFFX1 DFF_271_Q_reg ( .D(g28736), .SI(g423), .SE(test_se), .CLK(CK), .Q(
        test_so17), .QN() );
  SDFFX1 DFF_272_Q_reg ( .D(g28745), .SI(test_si18), .SE(test_se), .CLK(CK), 
        .Q(g428), .QN() );
  SDFFX1 DFF_273_Q_reg ( .D(g28754), .SI(g428), .SE(test_se), .CLK(CK), .Q(
        g426), .QN() );
  SDFFX1 DFF_274_Q_reg ( .D(g26803), .SI(g426), .SE(test_se), .CLK(CK), .Q(
        g429), .QN() );
  SDFFX1 DFF_275_Q_reg ( .D(g26804), .SI(g429), .SE(test_se), .CLK(CK), .Q(
        g432), .QN() );
  SDFFX1 DFF_276_Q_reg ( .D(g26807), .SI(g432), .SE(test_se), .CLK(CK), .Q(
        g435), .QN() );
  SDFFX1 DFF_277_Q_reg ( .D(g26805), .SI(g435), .SE(test_se), .CLK(CK), .Q(
        g438), .QN() );
  SDFFX1 DFF_278_Q_reg ( .D(g26808), .SI(g438), .SE(test_se), .CLK(CK), .Q(
        g441), .QN() );
  SDFFX1 DFF_279_Q_reg ( .D(g26812), .SI(g441), .SE(test_se), .CLK(CK), .Q(
        g444), .QN() );
  SDFFX1 DFF_280_Q_reg ( .D(g27759), .SI(g444), .SE(test_se), .CLK(CK), .Q(
        g448), .QN() );
  SDFFX1 DFF_281_Q_reg ( .D(g27760), .SI(g448), .SE(test_se), .CLK(CK), .Q(
        g449), .QN() );
  SDFFX1 DFF_282_Q_reg ( .D(g27762), .SI(g449), .SE(test_se), .CLK(CK), .Q(
        g447), .QN() );
  SDFFX1 DFF_283_Q_reg ( .D(g29606), .SI(g447), .SE(test_se), .CLK(CK), .Q(
        g312), .QN() );
  SDFFX1 DFF_284_Q_reg ( .D(g29608), .SI(g312), .SE(test_se), .CLK(CK), .Q(
        g313), .QN() );
  SDFFX1 DFF_285_Q_reg ( .D(g29611), .SI(g313), .SE(test_se), .CLK(CK), .Q(
        g314), .QN() );
  SDFFX1 DFF_286_Q_reg ( .D(g30699), .SI(g314), .SE(test_se), .CLK(CK), .Q(
        g315), .QN() );
  SDFFX1 DFF_287_Q_reg ( .D(g30700), .SI(g315), .SE(test_se), .CLK(CK), .Q(
        test_so18), .QN() );
  SDFFX1 DFF_288_Q_reg ( .D(g30702), .SI(test_si19), .SE(test_se), .CLK(CK), 
        .Q(g317), .QN() );
  SDFFX1 DFF_289_Q_reg ( .D(g30455), .SI(g317), .SE(test_se), .CLK(CK), .Q(
        g318), .QN() );
  SDFFX1 DFF_290_Q_reg ( .D(g30468), .SI(g318), .SE(test_se), .CLK(CK), .Q(
        g319), .QN() );
  SDFFX1 DFF_291_Q_reg ( .D(g30482), .SI(g319), .SE(test_se), .CLK(CK), .Q(
        g320), .QN() );
  SDFFX1 DFF_292_Q_reg ( .D(g29167), .SI(g320), .SE(test_se), .CLK(CK), .Q(
        g322), .QN() );
  SDFFX1 DFF_293_Q_reg ( .D(g29169), .SI(g322), .SE(test_se), .CLK(CK), .Q(
        g323), .QN() );
  SDFFX1 DFF_294_Q_reg ( .D(g29172), .SI(g323), .SE(test_se), .CLK(CK), .Q(
        g321), .QN() );
  SDFFX1 DFF_295_Q_reg ( .D(g26655), .SI(g321), .SE(test_se), .CLK(CK), .Q(
        g403), .QN() );
  SDFFX1 DFF_296_Q_reg ( .D(g26659), .SI(g403), .SE(test_se), .CLK(CK), .Q(
        g404), .QN() );
  SDFFX1 DFF_297_Q_reg ( .D(g26664), .SI(g404), .SE(test_se), .CLK(CK), .Q(
        g402), .QN() );
  SDFFX1 DFF_298_Q_reg ( .D(n4290), .SI(g402), .SE(test_se), .CLK(CK), .Q(g450), .QN() );
  SDFFX1 DFF_299_Q_reg ( .D(g450), .SI(g450), .SE(test_se), .CLK(CK), .Q(n8066), .QN(DFF_299_n1) );
  SDFFX1 DFF_300_Q_reg ( .D(n4569), .SI(n8066), .SE(test_se), .CLK(CK), .Q(
        g452), .QN() );
  SDFFX1 DFF_301_Q_reg ( .D(g452), .SI(g452), .SE(test_se), .CLK(CK), .Q(n8065), .QN(DFF_301_n1) );
  SDFFX1 DFF_302_Q_reg ( .D(n4561), .SI(n8065), .SE(test_se), .CLK(CK), .Q(
        g454), .QN() );
  SDFFX1 DFF_303_Q_reg ( .D(g454), .SI(g454), .SE(test_se), .CLK(CK), .Q(
        test_so19), .QN(DFF_303_n1) );
  SDFFX1 DFF_304_Q_reg ( .D(n4328), .SI(test_si20), .SE(test_se), .CLK(CK), 
        .Q(g280), .QN() );
  SDFFX1 DFF_305_Q_reg ( .D(g280), .SI(g280), .SE(test_se), .CLK(CK), .Q(n8062), .QN(DFF_305_n1) );
  SDFFX1 DFF_306_Q_reg ( .D(n4392), .SI(n8062), .SE(test_se), .CLK(CK), .Q(
        g282), .QN() );
  SDFFX1 DFF_307_Q_reg ( .D(g282), .SI(g282), .SE(test_se), .CLK(CK), .Q(n8061), .QN(DFF_307_n1) );
  SDFFX1 DFF_308_Q_reg ( .D(n4322), .SI(n8061), .SE(test_se), .CLK(CK), .Q(
        g284), .QN() );
  SDFFX1 DFF_309_Q_reg ( .D(g284), .SI(g284), .SE(test_se), .CLK(CK), .Q(n8060), .QN(DFF_309_n1) );
  SDFFX1 DFF_310_Q_reg ( .D(n4376), .SI(n8060), .SE(test_se), .CLK(CK), .Q(
        g286), .QN() );
  SDFFX1 DFF_311_Q_reg ( .D(g286), .SI(g286), .SE(test_se), .CLK(CK), .Q(n8059), .QN(DFF_311_n1) );
  SDFFX1 DFF_312_Q_reg ( .D(n4380), .SI(n8059), .SE(test_se), .CLK(CK), .Q(
        g288), .QN() );
  SDFFX1 DFF_313_Q_reg ( .D(g288), .SI(g288), .SE(test_se), .CLK(CK), .Q(n8058), .QN(DFF_313_n1) );
  SDFFX1 DFF_314_Q_reg ( .D(g2857), .SI(n8058), .SE(test_se), .CLK(CK), .Q(
        g290), .QN() );
  SDFFX1 DFF_315_Q_reg ( .D(g290), .SI(g290), .SE(test_se), .CLK(CK), .Q(n8057), .QN(n4485) );
  SDFFX1 DFF_316_Q_reg ( .D(n4282), .SI(n8057), .SE(test_se), .CLK(CK), .Q(
        n8056), .QN(n4430) );
  SDFFX1 DFF_317_Q_reg ( .D(g21346), .SI(n8056), .SE(test_se), .CLK(CK), .Q(
        g305), .QN() );
  SDFFX1 DFF_328_Q_reg ( .D(n4278), .SI(g305), .SE(test_se), .CLK(CK), .Q(
        n8055), .QN(DFF_328_n1) );
  SDFFX1 DFF_329_Q_reg ( .D(g354), .SI(n8055), .SE(test_se), .CLK(CK), .Q(
        test_so20), .QN() );
  SDFFX1 DFF_330_Q_reg ( .D(test_so20), .SI(test_si21), .SE(test_se), .CLK(CK), 
        .Q(g349), .QN() );
  SDFFX1 DFF_331_Q_reg ( .D(g343), .SI(g349), .SE(test_se), .CLK(CK), .Q(g350), 
        .QN() );
  SDFFX1 DFF_332_Q_reg ( .D(g350), .SI(g350), .SE(test_se), .CLK(CK), .Q(g351), 
        .QN() );
  SDFFX1 DFF_333_Q_reg ( .D(test_so16), .SI(g351), .SE(test_se), .CLK(CK), .Q(
        g352), .QN() );
  SDFFX1 DFF_334_Q_reg ( .D(g352), .SI(g352), .SE(test_se), .CLK(CK), .Q(g353), 
        .QN() );
  SDFFX1 DFF_335_Q_reg ( .D(g369), .SI(g353), .SE(test_se), .CLK(CK), .Q(g357), 
        .QN() );
  SDFFX1 DFF_336_Q_reg ( .D(g357), .SI(g357), .SE(test_se), .CLK(CK), .Q(g364), 
        .QN() );
  SDFFX1 DFF_337_Q_reg ( .D(g358), .SI(g364), .SE(test_se), .CLK(CK), .Q(g365), 
        .QN() );
  SDFFX1 DFF_338_Q_reg ( .D(g365), .SI(g365), .SE(test_se), .CLK(CK), .Q(g366), 
        .QN() );
  SDFFX1 DFF_339_Q_reg ( .D(g361), .SI(g366), .SE(test_se), .CLK(CK), .Q(g367), 
        .QN() );
  SDFFX1 DFF_340_Q_reg ( .D(g367), .SI(g367), .SE(test_se), .CLK(CK), .Q(g368), 
        .QN() );
  SDFFX1 DFF_341_Q_reg ( .D(g384), .SI(g368), .SE(test_se), .CLK(CK), .Q(g372), 
        .QN() );
  SDFFX1 DFF_342_Q_reg ( .D(g372), .SI(g372), .SE(test_se), .CLK(CK), .Q(g379), 
        .QN() );
  SDFFX1 DFF_343_Q_reg ( .D(g373), .SI(g379), .SE(test_se), .CLK(CK), .Q(g380), 
        .QN() );
  SDFFX1 DFF_344_Q_reg ( .D(g380), .SI(g380), .SE(test_se), .CLK(CK), .Q(g381), 
        .QN() );
  SDFFX1 DFF_345_Q_reg ( .D(g376), .SI(g381), .SE(test_se), .CLK(CK), .Q(
        test_so21), .QN() );
  SDFFX1 DFF_346_Q_reg ( .D(test_so21), .SI(test_si22), .SE(test_se), .CLK(CK), 
        .Q(g383), .QN() );
  SDFFX1 DFF_347_Q_reg ( .D(g398), .SI(g383), .SE(test_se), .CLK(CK), .Q(g387), 
        .QN() );
  SDFFX1 DFF_348_Q_reg ( .D(g387), .SI(g387), .SE(test_se), .CLK(CK), .Q(g394), 
        .QN() );
  SDFFX1 DFF_349_Q_reg ( .D(g388), .SI(g394), .SE(test_se), .CLK(CK), .Q(g395), 
        .QN() );
  SDFFX1 DFF_350_Q_reg ( .D(g395), .SI(g395), .SE(test_se), .CLK(CK), .Q(g396), 
        .QN() );
  SDFFX1 DFF_351_Q_reg ( .D(g391), .SI(g396), .SE(test_se), .CLK(CK), .Q(g397), 
        .QN() );
  SDFFX1 DFF_352_Q_reg ( .D(g397), .SI(g397), .SE(test_se), .CLK(CK), .Q(g324), 
        .QN() );
  SDFFX1 DFF_353_Q_reg ( .D(n4598), .SI(g324), .SE(test_se), .CLK(CK), .Q(
        g5629), .QN() );
  SDFFX1 DFF_354_Q_reg ( .D(g5629), .SI(g5629), .SE(test_se), .CLK(CK), .Q(
        g5648), .QN() );
  SDFFX1 DFF_355_Q_reg ( .D(g5648), .SI(g5648), .SE(test_se), .CLK(CK), .Q(
        g337), .QN() );
  SDFFX1 DFF_356_Q_reg ( .D(n4598), .SI(g337), .SE(test_se), .CLK(CK), .Q(g545), .QN(n4298) );
  SDFFX1 DFF_357_Q_reg ( .D(g6485), .SI(g545), .SE(test_se), .CLK(CK), .Q(g551), .QN(n4372) );
  SDFFX1 DFF_358_Q_reg ( .D(n4636), .SI(g551), .SE(test_se), .CLK(CK), .Q(g550), .QN(n4313) );
  SDFFX1 DFF_359_Q_reg ( .D(g21842), .SI(g550), .SE(test_se), .CLK(CK), .Q(
        g554), .QN() );
  SDFFX1 DFF_360_Q_reg ( .D(g18678), .SI(g554), .SE(test_se), .CLK(CK), .Q(
        g557), .QN(n4360) );
  SDFFX1 DFF_361_Q_reg ( .D(g18726), .SI(g557), .SE(test_se), .CLK(CK), .Q(
        test_so22), .QN(n4310) );
  SDFFX1 DFF_362_Q_reg ( .D(g12487), .SI(test_si23), .SE(test_se), .CLK(CK), 
        .Q(g513), .QN() );
  SDFFX1 DFF_363_Q_reg ( .D(g513), .SI(g513), .SE(test_se), .CLK(CK), .Q(g523), 
        .QN() );
  SDFFX1 DFF_364_Q_reg ( .D(g523), .SI(g523), .SE(test_se), .CLK(CK), .Q(g524), 
        .QN() );
  SDFFX1 DFF_365_Q_reg ( .D(g455), .SI(g524), .SE(test_se), .CLK(CK), .Q(g564), 
        .QN() );
  SDFFX1 DFF_366_Q_reg ( .D(g564), .SI(g564), .SE(test_se), .CLK(CK), .Q(g569), 
        .QN() );
  SDFFX1 DFF_367_Q_reg ( .D(g458), .SI(g569), .SE(test_se), .CLK(CK), .Q(g570), 
        .QN() );
  SDFFX1 DFF_368_Q_reg ( .D(g570), .SI(g570), .SE(test_se), .CLK(CK), .Q(g571), 
        .QN() );
  SDFFX1 DFF_369_Q_reg ( .D(g461), .SI(g571), .SE(test_se), .CLK(CK), .Q(g572), 
        .QN() );
  SDFFX1 DFF_370_Q_reg ( .D(g572), .SI(g572), .SE(test_se), .CLK(CK), .Q(g573), 
        .QN() );
  SDFFX1 DFF_371_Q_reg ( .D(g465), .SI(g573), .SE(test_se), .CLK(CK), .Q(g574), 
        .QN() );
  SDFFX1 DFF_372_Q_reg ( .D(g574), .SI(g574), .SE(test_se), .CLK(CK), .Q(g565), 
        .QN() );
  SDFFX1 DFF_373_Q_reg ( .D(test_so24), .SI(g565), .SE(test_se), .CLK(CK), .Q(
        g566), .QN() );
  SDFFX1 DFF_374_Q_reg ( .D(g566), .SI(g566), .SE(test_se), .CLK(CK), .Q(g567), 
        .QN() );
  SDFFX1 DFF_375_Q_reg ( .D(g471), .SI(g567), .SE(test_se), .CLK(CK), .Q(g568), 
        .QN() );
  SDFFX1 DFF_376_Q_reg ( .D(g568), .SI(g568), .SE(test_se), .CLK(CK), .Q(g489), 
        .QN() );
  SDFFX1 DFF_377_Q_reg ( .D(n4650), .SI(g489), .SE(test_se), .CLK(CK), .Q(
        g7909), .QN(n4462) );
  SDFFX1 DFF_378_Q_reg ( .D(g7909), .SI(test_si24), .SE(test_se), .CLK(CK), 
        .Q(g7956), .QN(n4461) );
  SDFFX1 DFF_379_Q_reg ( .D(g7956), .SI(g7956), .SE(test_se), .CLK(CK), .Q(
        g485), .QN(n4466) );
  SDFFX1 DFF_380_Q_reg ( .D(g23067), .SI(g485), .SE(test_se), .CLK(CK), .Q(
        g486), .QN() );
  SDFFX1 DFF_381_Q_reg ( .D(g23093), .SI(g486), .SE(test_se), .CLK(CK), .Q(
        g487), .QN() );
  SDFFX1 DFF_382_Q_reg ( .D(g23117), .SI(g487), .SE(test_se), .CLK(CK), .Q(
        g488), .QN() );
  SDFFX1 DFF_383_Q_reg ( .D(g23385), .SI(g488), .SE(test_se), .CLK(CK), .Q(
        g455), .QN() );
  SDFFX1 DFF_384_Q_reg ( .D(g23399), .SI(g455), .SE(test_se), .CLK(CK), .Q(
        g458), .QN() );
  SDFFX1 DFF_385_Q_reg ( .D(g24174), .SI(g458), .SE(test_se), .CLK(CK), .Q(
        g461), .QN() );
  SDFFX1 DFF_386_Q_reg ( .D(g24178), .SI(g461), .SE(test_se), .CLK(CK), .Q(
        g477), .QN() );
  SDFFX1 DFF_387_Q_reg ( .D(g24207), .SI(g477), .SE(test_se), .CLK(CK), .Q(
        g478), .QN() );
  SDFFX1 DFF_388_Q_reg ( .D(g24216), .SI(g478), .SE(test_se), .CLK(CK), .Q(
        g479), .QN() );
  SDFFX1 DFF_389_Q_reg ( .D(g23092), .SI(g479), .SE(test_se), .CLK(CK), .Q(
        g480), .QN() );
  SDFFX1 DFF_390_Q_reg ( .D(g23000), .SI(g480), .SE(test_se), .CLK(CK), .Q(
        g484), .QN() );
  SDFFX1 DFF_391_Q_reg ( .D(g23022), .SI(g484), .SE(test_se), .CLK(CK), .Q(
        g464), .QN() );
  SDFFX1 DFF_392_Q_reg ( .D(g24206), .SI(g464), .SE(test_se), .CLK(CK), .Q(
        g465), .QN() );
  SDFFX1 DFF_393_Q_reg ( .D(g24215), .SI(g465), .SE(test_se), .CLK(CK), .Q(
        test_so24), .QN() );
  SDFFX1 DFF_394_Q_reg ( .D(g24228), .SI(test_si25), .SE(test_se), .CLK(CK), 
        .Q(g471), .QN() );
  SDFFX1 DFF_395_Q_reg ( .D(g12457), .SI(g471), .SE(test_se), .CLK(CK), .Q(
        g528), .QN() );
  SDFFX1 DFF_396_Q_reg ( .D(g528), .SI(g528), .SE(test_se), .CLK(CK), .Q(g535), 
        .QN() );
  SDFFX1 DFF_397_Q_reg ( .D(g535), .SI(g535), .SE(test_se), .CLK(CK), .Q(g542), 
        .QN() );
  SDFFX1 DFF_398_Q_reg ( .D(g13149), .SI(g542), .SE(test_se), .CLK(CK), .Q(
        g543), .QN() );
  SDFFX1 DFF_399_Q_reg ( .D(g543), .SI(g543), .SE(test_se), .CLK(CK), .Q(g544), 
        .QN() );
  SDFFX1 DFF_400_Q_reg ( .D(g21851), .SI(g544), .SE(test_se), .CLK(CK), .Q(
        g548), .QN() );
  SDFFX1 DFF_401_Q_reg ( .D(g13111), .SI(g548), .SE(test_se), .CLK(CK), .Q(
        g549), .QN() );
  SDFFX1 DFF_402_Q_reg ( .D(g549), .SI(g549), .SE(test_se), .CLK(CK), .Q(g499), 
        .QN(n4541) );
  SDFFX1 DFF_403_Q_reg ( .D(g13160), .SI(g499), .SE(test_se), .CLK(CK), .Q(
        g558), .QN() );
  SDFFX1 DFF_404_Q_reg ( .D(g558), .SI(g558), .SE(test_se), .CLK(CK), .Q(g559), 
        .QN() );
  SDFFX1 DFF_405_Q_reg ( .D(g27261), .SI(g559), .SE(test_se), .CLK(CK), .Q(
        g576), .QN() );
  SDFFX1 DFF_406_Q_reg ( .D(g27268), .SI(g576), .SE(test_se), .CLK(CK), .Q(
        g577), .QN() );
  SDFFX1 DFF_407_Q_reg ( .D(g27279), .SI(g577), .SE(test_se), .CLK(CK), .Q(
        g575), .QN() );
  SDFFX1 DFF_408_Q_reg ( .D(g27269), .SI(g575), .SE(test_se), .CLK(CK), .Q(
        g579), .QN() );
  SDFFX1 DFF_409_Q_reg ( .D(g27280), .SI(g579), .SE(test_se), .CLK(CK), .Q(
        test_so25), .QN() );
  SDFFX1 DFF_410_Q_reg ( .D(g27294), .SI(test_si26), .SE(test_se), .CLK(CK), 
        .Q(g578), .QN() );
  SDFFX1 DFF_411_Q_reg ( .D(g27281), .SI(g578), .SE(test_se), .CLK(CK), .Q(
        g582), .QN() );
  SDFFX1 DFF_412_Q_reg ( .D(g27295), .SI(g582), .SE(test_se), .CLK(CK), .Q(
        g583), .QN() );
  SDFFX1 DFF_413_Q_reg ( .D(g27311), .SI(g583), .SE(test_se), .CLK(CK), .Q(
        g581), .QN() );
  SDFFX1 DFF_414_Q_reg ( .D(g27296), .SI(g581), .SE(test_se), .CLK(CK), .Q(
        g585), .QN() );
  SDFFX1 DFF_415_Q_reg ( .D(g27312), .SI(g585), .SE(test_se), .CLK(CK), .Q(
        g586), .QN() );
  SDFFX1 DFF_416_Q_reg ( .D(g27327), .SI(g586), .SE(test_se), .CLK(CK), .Q(
        g584), .QN() );
  SDFFX1 DFF_417_Q_reg ( .D(g24491), .SI(g584), .SE(test_se), .CLK(CK), .Q(
        g587), .QN() );
  SDFFX1 DFF_418_Q_reg ( .D(g24498), .SI(g587), .SE(test_se), .CLK(CK), .Q(
        g590), .QN() );
  SDFFX1 DFF_419_Q_reg ( .D(g24507), .SI(g590), .SE(test_se), .CLK(CK), .Q(
        g593), .QN() );
  SDFFX1 DFF_420_Q_reg ( .D(g24499), .SI(g593), .SE(test_se), .CLK(CK), .Q(
        g596), .QN() );
  SDFFX1 DFF_421_Q_reg ( .D(g24508), .SI(g596), .SE(test_se), .CLK(CK), .Q(
        g599), .QN() );
  SDFFX1 DFF_422_Q_reg ( .D(g24519), .SI(g599), .SE(test_se), .CLK(CK), .Q(
        g602), .QN() );
  SDFFX1 DFF_423_Q_reg ( .D(g28345), .SI(g602), .SE(test_se), .CLK(CK), .Q(
        g614), .QN() );
  SDFFX1 DFF_424_Q_reg ( .D(g28349), .SI(g614), .SE(test_se), .CLK(CK), .Q(
        g617), .QN() );
  SDFFX1 DFF_425_Q_reg ( .D(g28353), .SI(g617), .SE(test_se), .CLK(CK), .Q(
        test_so26), .QN() );
  SDFFX1 DFF_426_Q_reg ( .D(g28342), .SI(test_si27), .SE(test_se), .CLK(CK), 
        .Q(g605), .QN() );
  SDFFX1 DFF_427_Q_reg ( .D(g28344), .SI(g605), .SE(test_se), .CLK(CK), .Q(
        g608), .QN() );
  SDFFX1 DFF_428_Q_reg ( .D(g28348), .SI(g608), .SE(test_se), .CLK(CK), .Q(
        g611), .QN() );
  SDFFX1 DFF_429_Q_reg ( .D(g26541), .SI(g611), .SE(test_se), .CLK(CK), .Q(
        g490), .QN() );
  SDFFX1 DFF_430_Q_reg ( .D(g26545), .SI(g490), .SE(test_se), .CLK(CK), .Q(
        g493), .QN() );
  SDFFX1 DFF_431_Q_reg ( .D(g26553), .SI(g493), .SE(test_se), .CLK(CK), .Q(
        g496), .QN() );
  SDFFX1 DFF_432_Q_reg ( .D(g499), .SI(g496), .SE(test_se), .CLK(CK), .Q(g506), 
        .QN(n4570) );
  SDFFX1 DFF_433_Q_reg ( .D(g22578), .SI(g506), .SE(test_se), .CLK(CK), .Q(
        n4571), .QN() );
  SDFFX1 DFF_442_Q_reg ( .D(n1828), .SI(n4571), .SE(test_se), .CLK(CK), .Q(
        g16297), .QN() );
  SDFFX1 DFF_443_Q_reg ( .D(g16297), .SI(g16297), .SE(test_se), .CLK(CK), .Q(
        g525), .QN() );
  SDFFX1 DFF_444_Q_reg ( .D(DFF_299_n1), .SI(g525), .SE(test_se), .CLK(CK), 
        .Q(n8047), .QN(DFF_444_n1) );
  SDFFX1 DFF_445_Q_reg ( .D(DFF_301_n1), .SI(n8047), .SE(test_se), .CLK(CK), 
        .Q(n8046), .QN(DFF_445_n1) );
  SDFFX1 DFF_446_Q_reg ( .D(DFF_303_n1), .SI(n8046), .SE(test_se), .CLK(CK), 
        .Q(n8045), .QN(DFF_446_n1) );
  SDFFX1 DFF_447_Q_reg ( .D(DFF_305_n1), .SI(n8045), .SE(test_se), .CLK(CK), 
        .Q(n8044), .QN(DFF_447_n1) );
  SDFFX1 DFF_448_Q_reg ( .D(DFF_307_n1), .SI(n8044), .SE(test_se), .CLK(CK), 
        .Q(n8043), .QN(DFF_448_n1) );
  SDFFX1 DFF_449_Q_reg ( .D(DFF_309_n1), .SI(n8043), .SE(test_se), .CLK(CK), 
        .Q(test_so27), .QN(DFF_449_n1) );
  SDFFX1 DFF_450_Q_reg ( .D(DFF_311_n1), .SI(test_si28), .SE(test_se), .CLK(CK), .Q(g536), .QN() );
  SDFFX1 DFF_451_Q_reg ( .D(DFF_313_n1), .SI(g536), .SE(test_se), .CLK(CK), 
        .Q(g537), .QN() );
  SDFFX1 DFF_452_Q_reg ( .D(g24059), .SI(g537), .SE(test_se), .CLK(CK), .Q(
        g538), .QN(n4492) );
  SDFFX1 DFF_453_Q_reg ( .D(n4485), .SI(g538), .SE(test_se), .CLK(CK), .Q(
        n8040), .QN(DFF_453_n1) );
  SDFFX1 DFF_455_Q_reg ( .D(g6677), .SI(g6677), .SE(test_se), .CLK(CK), .Q(
        g6911), .QN(n4359) );
  SDFFX1 DFF_456_Q_reg ( .D(g6911), .SI(g6911), .SE(test_se), .CLK(CK), .Q(
        g629), .QN(n4295) );
  SDFFX1 DFF_457_Q_reg ( .D(g16654), .SI(g629), .SE(test_se), .CLK(CK), .Q(
        g630), .QN() );
  SDFFX1 DFF_458_Q_reg ( .D(g20314), .SI(g630), .SE(test_se), .CLK(CK), .Q(
        g659), .QN(n4429) );
  SDFFX1 DFF_459_Q_reg ( .D(g20682), .SI(g659), .SE(test_se), .CLK(CK), .Q(
        g640), .QN(n4404) );
  SDFFX1 DFF_460_Q_reg ( .D(g23136), .SI(g640), .SE(test_se), .CLK(CK), .Q(
        g633), .QN(n4478) );
  SDFFX1 DFF_461_Q_reg ( .D(g23324), .SI(g633), .SE(test_se), .CLK(CK), .Q(
        g653), .QN(n4422) );
  SDFFX1 DFF_462_Q_reg ( .D(g24426), .SI(g653), .SE(test_se), .CLK(CK), .Q(
        g646), .QN(n4414) );
  SDFFX1 DFF_463_Q_reg ( .D(g25185), .SI(g646), .SE(test_se), .CLK(CK), .Q(
        g660), .QN(n4403) );
  SDFFX1 DFF_464_Q_reg ( .D(g26660), .SI(g660), .SE(test_se), .CLK(CK), .Q(
        g672), .QN(n4413) );
  SDFFX1 DFF_465_Q_reg ( .D(g26776), .SI(g672), .SE(test_se), .CLK(CK), .Q(
        test_so28), .QN(n4470) );
  SDFFX1 DFF_466_Q_reg ( .D(g27672), .SI(test_si29), .SE(test_se), .CLK(CK), 
        .Q(g679), .QN(n4477) );
  SDFFX1 DFF_467_Q_reg ( .D(g28199), .SI(g679), .SE(test_se), .CLK(CK), .Q(
        g686), .QN(n4396) );
  SDFFX1 DFF_468_Q_reg ( .D(g28668), .SI(g686), .SE(test_se), .CLK(CK), .Q(
        g692), .QN(n4418) );
  SDFFX1 DFF_469_Q_reg ( .D(g20875), .SI(g692), .SE(test_se), .CLK(CK), .Q(
        g699), .QN() );
  SDFFX1 DFF_470_Q_reg ( .D(g20879), .SI(g699), .SE(test_se), .CLK(CK), .Q(
        g700), .QN() );
  SDFFX1 DFF_471_Q_reg ( .D(g20891), .SI(g700), .SE(test_se), .CLK(CK), .Q(
        g698), .QN() );
  SDFFX1 DFF_472_Q_reg ( .D(g20880), .SI(g698), .SE(test_se), .CLK(CK), .Q(
        g702), .QN() );
  SDFFX1 DFF_473_Q_reg ( .D(g20892), .SI(g702), .SE(test_se), .CLK(CK), .Q(
        g703), .QN() );
  SDFFX1 DFF_474_Q_reg ( .D(g20901), .SI(g703), .SE(test_se), .CLK(CK), .Q(
        g701), .QN() );
  SDFFX1 DFF_475_Q_reg ( .D(g20893), .SI(g701), .SE(test_se), .CLK(CK), .Q(
        g705), .QN() );
  SDFFX1 DFF_476_Q_reg ( .D(g20902), .SI(g705), .SE(test_se), .CLK(CK), .Q(
        g706), .QN() );
  SDFFX1 DFF_477_Q_reg ( .D(g20921), .SI(g706), .SE(test_se), .CLK(CK), .Q(
        g704), .QN() );
  SDFFX1 DFF_478_Q_reg ( .D(g20903), .SI(g704), .SE(test_se), .CLK(CK), .Q(
        g708), .QN() );
  SDFFX1 DFF_479_Q_reg ( .D(g20922), .SI(g708), .SE(test_se), .CLK(CK), .Q(
        g709), .QN() );
  SDFFX1 DFF_480_Q_reg ( .D(g20944), .SI(g709), .SE(test_se), .CLK(CK), .Q(
        g707), .QN() );
  SDFFX1 DFF_481_Q_reg ( .D(g20923), .SI(g707), .SE(test_se), .CLK(CK), .Q(
        test_so29), .QN() );
  SDFFX1 DFF_482_Q_reg ( .D(g20945), .SI(test_si30), .SE(test_se), .CLK(CK), 
        .Q(g712), .QN() );
  SDFFX1 DFF_483_Q_reg ( .D(g20966), .SI(g712), .SE(test_se), .CLK(CK), .Q(
        g710), .QN() );
  SDFFX1 DFF_484_Q_reg ( .D(g20946), .SI(g710), .SE(test_se), .CLK(CK), .Q(
        g714), .QN() );
  SDFFX1 DFF_485_Q_reg ( .D(g20967), .SI(g714), .SE(test_se), .CLK(CK), .Q(
        g715), .QN() );
  SDFFX1 DFF_486_Q_reg ( .D(g20989), .SI(g715), .SE(test_se), .CLK(CK), .Q(
        g713), .QN() );
  SDFFX1 DFF_487_Q_reg ( .D(g20968), .SI(g713), .SE(test_se), .CLK(CK), .Q(
        g717), .QN() );
  SDFFX1 DFF_488_Q_reg ( .D(g20990), .SI(g717), .SE(test_se), .CLK(CK), .Q(
        g718), .QN() );
  SDFFX1 DFF_489_Q_reg ( .D(g21009), .SI(g718), .SE(test_se), .CLK(CK), .Q(
        g716), .QN() );
  SDFFX1 DFF_490_Q_reg ( .D(g20991), .SI(g716), .SE(test_se), .CLK(CK), .Q(
        g720), .QN() );
  SDFFX1 DFF_491_Q_reg ( .D(g21010), .SI(g720), .SE(test_se), .CLK(CK), .Q(
        g721), .QN() );
  SDFFX1 DFF_492_Q_reg ( .D(g21031), .SI(g721), .SE(test_se), .CLK(CK), .Q(
        g719), .QN() );
  SDFFX1 DFF_493_Q_reg ( .D(g21011), .SI(g719), .SE(test_se), .CLK(CK), .Q(
        g723), .QN() );
  SDFFX1 DFF_494_Q_reg ( .D(g21032), .SI(g723), .SE(test_se), .CLK(CK), .Q(
        g724), .QN() );
  SDFFX1 DFF_495_Q_reg ( .D(g21051), .SI(g724), .SE(test_se), .CLK(CK), .Q(
        g722), .QN() );
  SDFFX1 DFF_496_Q_reg ( .D(g20876), .SI(g722), .SE(test_se), .CLK(CK), .Q(
        g726), .QN() );
  SDFFX1 DFF_497_Q_reg ( .D(g20881), .SI(g726), .SE(test_se), .CLK(CK), .Q(
        test_so30), .QN() );
  SDFFX1 DFF_498_Q_reg ( .D(g20894), .SI(test_si31), .SE(test_se), .CLK(CK), 
        .Q(g725), .QN() );
  SDFFX1 DFF_499_Q_reg ( .D(g20924), .SI(g725), .SE(test_se), .CLK(CK), .Q(
        g729), .QN() );
  SDFFX1 DFF_500_Q_reg ( .D(g20947), .SI(g729), .SE(test_se), .CLK(CK), .Q(
        g730), .QN() );
  SDFFX1 DFF_501_Q_reg ( .D(g20969), .SI(g730), .SE(test_se), .CLK(CK), .Q(
        g728), .QN() );
  SDFFX1 DFF_502_Q_reg ( .D(g20948), .SI(g728), .SE(test_se), .CLK(CK), .Q(
        g732), .QN() );
  SDFFX1 DFF_503_Q_reg ( .D(g20970), .SI(g732), .SE(test_se), .CLK(CK), .Q(
        g733), .QN() );
  SDFFX1 DFF_504_Q_reg ( .D(g20992), .SI(g733), .SE(test_se), .CLK(CK), .Q(
        g731), .QN() );
  SDFFX1 DFF_505_Q_reg ( .D(g25260), .SI(g731), .SE(test_se), .CLK(CK), .Q(
        g735), .QN() );
  SDFFX1 DFF_506_Q_reg ( .D(g25262), .SI(g735), .SE(test_se), .CLK(CK), .Q(
        g736), .QN() );
  SDFFX1 DFF_507_Q_reg ( .D(g25266), .SI(g736), .SE(test_se), .CLK(CK), .Q(
        g734), .QN() );
  SDFFX1 DFF_508_Q_reg ( .D(g22218), .SI(g734), .SE(test_se), .CLK(CK), .Q(
        g738), .QN() );
  SDFFX1 DFF_509_Q_reg ( .D(g22231), .SI(g738), .SE(test_se), .CLK(CK), .Q(
        g739), .QN() );
  SDFFX1 DFF_510_Q_reg ( .D(g22242), .SI(g739), .SE(test_se), .CLK(CK), .Q(
        g737), .QN() );
  SDFFX1 DFF_511_Q_reg ( .D(n4650), .SI(g737), .SE(test_se), .CLK(CK), .Q(
        g6368), .QN(n4323) );
  SDFFX1 DFF_512_Q_reg ( .D(n4592), .SI(g6368), .SE(test_se), .CLK(CK), .Q(
        g6518), .QN(n4312) );
  SDFFX1 DFF_513_Q_reg ( .D(n4591), .SI(g6518), .SE(test_se), .CLK(CK), .Q(
        test_so31), .QN(n4362) );
  SDFFX1 DFF_514_Q_reg ( .D(g22126), .SI(test_si32), .SE(test_se), .CLK(CK), 
        .Q(g818), .QN() );
  SDFFX1 DFF_515_Q_reg ( .D(g22145), .SI(g818), .SE(test_se), .CLK(CK), .Q(
        g819), .QN() );
  SDFFX1 DFF_516_Q_reg ( .D(g22162), .SI(g819), .SE(test_se), .CLK(CK), .Q(
        g817), .QN() );
  SDFFX1 DFF_517_Q_reg ( .D(g22146), .SI(g817), .SE(test_se), .CLK(CK), .Q(
        g821), .QN() );
  SDFFX1 DFF_518_Q_reg ( .D(g22163), .SI(g821), .SE(test_se), .CLK(CK), .Q(
        g822), .QN() );
  SDFFX1 DFF_519_Q_reg ( .D(g22177), .SI(g822), .SE(test_se), .CLK(CK), .Q(
        g820), .QN() );
  SDFFX1 DFF_520_Q_reg ( .D(g22029), .SI(g820), .SE(test_se), .CLK(CK), .Q(
        g830), .QN() );
  SDFFX1 DFF_521_Q_reg ( .D(g22033), .SI(g830), .SE(test_se), .CLK(CK), .Q(
        g831), .QN() );
  SDFFX1 DFF_522_Q_reg ( .D(g22040), .SI(g831), .SE(test_se), .CLK(CK), .Q(
        g829), .QN() );
  SDFFX1 DFF_523_Q_reg ( .D(g22034), .SI(g829), .SE(test_se), .CLK(CK), .Q(
        g833), .QN() );
  SDFFX1 DFF_524_Q_reg ( .D(g22041), .SI(g833), .SE(test_se), .CLK(CK), .Q(
        g834), .QN() );
  SDFFX1 DFF_525_Q_reg ( .D(g22054), .SI(g834), .SE(test_se), .CLK(CK), .Q(
        g832), .QN() );
  SDFFX1 DFF_526_Q_reg ( .D(g22042), .SI(g832), .SE(test_se), .CLK(CK), .Q(
        g836), .QN() );
  SDFFX1 DFF_527_Q_reg ( .D(g22055), .SI(g836), .SE(test_se), .CLK(CK), .Q(
        g837), .QN() );
  SDFFX1 DFF_528_Q_reg ( .D(g22066), .SI(g837), .SE(test_se), .CLK(CK), .Q(
        g835), .QN() );
  SDFFX1 DFF_529_Q_reg ( .D(g22056), .SI(g835), .SE(test_se), .CLK(CK), .Q(
        test_so32), .QN() );
  SDFFX1 DFF_530_Q_reg ( .D(g22067), .SI(test_si33), .SE(test_se), .CLK(CK), 
        .Q(g840), .QN() );
  SDFFX1 DFF_531_Q_reg ( .D(g22087), .SI(g840), .SE(test_se), .CLK(CK), .Q(
        g838), .QN() );
  SDFFX1 DFF_532_Q_reg ( .D(g22068), .SI(g838), .SE(test_se), .CLK(CK), .Q(
        g842), .QN() );
  SDFFX1 DFF_533_Q_reg ( .D(g22088), .SI(g842), .SE(test_se), .CLK(CK), .Q(
        g843), .QN() );
  SDFFX1 DFF_534_Q_reg ( .D(g22104), .SI(g843), .SE(test_se), .CLK(CK), .Q(
        g841), .QN() );
  SDFFX1 DFF_535_Q_reg ( .D(g22089), .SI(g841), .SE(test_se), .CLK(CK), .Q(
        g845), .QN() );
  SDFFX1 DFF_536_Q_reg ( .D(g22105), .SI(g845), .SE(test_se), .CLK(CK), .Q(
        g846), .QN() );
  SDFFX1 DFF_537_Q_reg ( .D(g22127), .SI(g846), .SE(test_se), .CLK(CK), .Q(
        g844), .QN() );
  SDFFX1 DFF_538_Q_reg ( .D(g22106), .SI(g844), .SE(test_se), .CLK(CK), .Q(
        g848), .QN() );
  SDFFX1 DFF_539_Q_reg ( .D(g22128), .SI(g848), .SE(test_se), .CLK(CK), .Q(
        g849), .QN() );
  SDFFX1 DFF_540_Q_reg ( .D(g22147), .SI(g849), .SE(test_se), .CLK(CK), .Q(
        g847), .QN() );
  SDFFX1 DFF_541_Q_reg ( .D(g22129), .SI(g847), .SE(test_se), .CLK(CK), .Q(
        g851), .QN() );
  SDFFX1 DFF_542_Q_reg ( .D(g22148), .SI(g851), .SE(test_se), .CLK(CK), .Q(
        g852), .QN() );
  SDFFX1 DFF_543_Q_reg ( .D(g22164), .SI(g852), .SE(test_se), .CLK(CK), .Q(
        g850), .QN() );
  SDFFX1 DFF_544_Q_reg ( .D(g25209), .SI(g850), .SE(test_se), .CLK(CK), .Q(
        g857), .QN() );
  SDFFX1 DFF_545_Q_reg ( .D(g25214), .SI(g857), .SE(test_se), .CLK(CK), .Q(
        test_so33), .QN() );
  SDFFX1 DFF_546_Q_reg ( .D(g25221), .SI(test_si34), .SE(test_se), .CLK(CK), 
        .Q(g856), .QN() );
  SDFFX1 DFF_547_Q_reg ( .D(g25215), .SI(g856), .SE(test_se), .CLK(CK), .Q(
        g860), .QN() );
  SDFFX1 DFF_548_Q_reg ( .D(g25222), .SI(g860), .SE(test_se), .CLK(CK), .Q(
        g861), .QN() );
  SDFFX1 DFF_549_Q_reg ( .D(g25230), .SI(g861), .SE(test_se), .CLK(CK), .Q(
        g859), .QN() );
  SDFFX1 DFF_550_Q_reg ( .D(g25223), .SI(g859), .SE(test_se), .CLK(CK), .Q(
        g863), .QN() );
  SDFFX1 DFF_551_Q_reg ( .D(g25231), .SI(g863), .SE(test_se), .CLK(CK), .Q(
        g864), .QN() );
  SDFFX1 DFF_552_Q_reg ( .D(g25240), .SI(g864), .SE(test_se), .CLK(CK), .Q(
        g862), .QN() );
  SDFFX1 DFF_553_Q_reg ( .D(g25232), .SI(g862), .SE(test_se), .CLK(CK), .Q(
        g866), .QN() );
  SDFFX1 DFF_554_Q_reg ( .D(g25241), .SI(g866), .SE(test_se), .CLK(CK), .Q(
        g867), .QN() );
  SDFFX1 DFF_555_Q_reg ( .D(g25248), .SI(g867), .SE(test_se), .CLK(CK), .Q(
        g865), .QN() );
  SDFFX1 DFF_556_Q_reg ( .D(g30269), .SI(g865), .SE(test_se), .CLK(CK), .Q(
        g873), .QN() );
  SDFFX1 DFF_557_Q_reg ( .D(g30277), .SI(g873), .SE(test_se), .CLK(CK), .Q(
        g876), .QN() );
  SDFFX1 DFF_558_Q_reg ( .D(g30285), .SI(g876), .SE(test_se), .CLK(CK), .Q(
        g879), .QN() );
  SDFFX1 DFF_559_Q_reg ( .D(g30643), .SI(g879), .SE(test_se), .CLK(CK), .Q(
        g918), .QN() );
  SDFFX1 DFF_560_Q_reg ( .D(g30648), .SI(g918), .SE(test_se), .CLK(CK), .Q(
        g921), .QN() );
  SDFFX1 DFF_561_Q_reg ( .D(g30654), .SI(g921), .SE(test_se), .CLK(CK), .Q(
        test_so34), .QN() );
  SDFFX1 DFF_562_Q_reg ( .D(g30676), .SI(test_si35), .SE(test_se), .CLK(CK), 
        .Q(g882), .QN() );
  SDFFX1 DFF_563_Q_reg ( .D(g30681), .SI(g882), .SE(test_se), .CLK(CK), .Q(
        g885), .QN() );
  SDFFX1 DFF_564_Q_reg ( .D(g30687), .SI(g885), .SE(test_se), .CLK(CK), .Q(
        g888), .QN() );
  SDFFX1 DFF_565_Q_reg ( .D(g30649), .SI(g888), .SE(test_se), .CLK(CK), .Q(
        g927), .QN() );
  SDFFX1 DFF_566_Q_reg ( .D(g30655), .SI(g927), .SE(test_se), .CLK(CK), .Q(
        g930), .QN() );
  SDFFX1 DFF_567_Q_reg ( .D(g30662), .SI(g930), .SE(test_se), .CLK(CK), .Q(
        g933), .QN() );
  SDFFX1 DFF_568_Q_reg ( .D(g30286), .SI(g933), .SE(test_se), .CLK(CK), .Q(
        g891), .QN() );
  SDFFX1 DFF_569_Q_reg ( .D(g30293), .SI(g891), .SE(test_se), .CLK(CK), .Q(
        g894), .QN() );
  SDFFX1 DFF_570_Q_reg ( .D(g30298), .SI(g894), .SE(test_se), .CLK(CK), .Q(
        g897), .QN() );
  SDFFX1 DFF_571_Q_reg ( .D(g30259), .SI(g897), .SE(test_se), .CLK(CK), .Q(
        g936), .QN() );
  SDFFX1 DFF_572_Q_reg ( .D(g30264), .SI(g936), .SE(test_se), .CLK(CK), .Q(
        g939), .QN() );
  SDFFX1 DFF_573_Q_reg ( .D(g30270), .SI(g939), .SE(test_se), .CLK(CK), .Q(
        g942), .QN() );
  SDFFX1 DFF_574_Q_reg ( .D(g30247), .SI(g942), .SE(test_se), .CLK(CK), .Q(
        g900), .QN() );
  SDFFX1 DFF_575_Q_reg ( .D(g30249), .SI(g900), .SE(test_se), .CLK(CK), .Q(
        g903), .QN() );
  SDFFX1 DFF_576_Q_reg ( .D(g30251), .SI(g903), .SE(test_se), .CLK(CK), .Q(
        g906), .QN() );
  SDFFX1 DFF_577_Q_reg ( .D(g30265), .SI(g906), .SE(test_se), .CLK(CK), .Q(
        test_so35), .QN() );
  SDFFX1 DFF_578_Q_reg ( .D(g30271), .SI(test_si36), .SE(test_se), .CLK(CK), 
        .Q(g948), .QN() );
  SDFFX1 DFF_579_Q_reg ( .D(g30278), .SI(g948), .SE(test_se), .CLK(CK), .Q(
        g951), .QN() );
  SDFFX1 DFF_580_Q_reg ( .D(g30638), .SI(g951), .SE(test_se), .CLK(CK), .Q(
        g909), .QN() );
  SDFFX1 DFF_581_Q_reg ( .D(g30642), .SI(g909), .SE(test_se), .CLK(CK), .Q(
        g912), .QN() );
  SDFFX1 DFF_582_Q_reg ( .D(g30647), .SI(g912), .SE(test_se), .CLK(CK), .Q(
        g915), .QN() );
  SDFFX1 DFF_583_Q_reg ( .D(g30670), .SI(g915), .SE(test_se), .CLK(CK), .Q(
        g954), .QN() );
  SDFFX1 DFF_584_Q_reg ( .D(g30677), .SI(g954), .SE(test_se), .CLK(CK), .Q(
        g957), .QN() );
  SDFFX1 DFF_585_Q_reg ( .D(g30682), .SI(g957), .SE(test_se), .CLK(CK), .Q(
        g960), .QN() );
  SDFFX1 DFF_586_Q_reg ( .D(g25042), .SI(g960), .SE(test_se), .CLK(CK), .Q(
        g780), .QN() );
  SDFFX1 DFF_587_Q_reg ( .D(g25935), .SI(g780), .SE(test_se), .CLK(CK), .Q(
        g776), .QN() );
  SDFFX1 DFF_588_Q_reg ( .D(g26530), .SI(g776), .SE(test_se), .CLK(CK), .Q(
        g771), .QN() );
  SDFFX1 DFF_589_Q_reg ( .D(g27123), .SI(g771), .SE(test_se), .CLK(CK), .Q(
        g767), .QN() );
  SDFFX1 DFF_590_Q_reg ( .D(g27603), .SI(g767), .SE(test_se), .CLK(CK), .Q(
        g762), .QN() );
  SDFFX1 DFF_591_Q_reg ( .D(g28146), .SI(g762), .SE(test_se), .CLK(CK), .Q(
        g758), .QN() );
  SDFFX1 DFF_592_Q_reg ( .D(g28635), .SI(g758), .SE(test_se), .CLK(CK), .Q(
        g753), .QN() );
  SDFFX1 DFF_593_Q_reg ( .D(g29110), .SI(g753), .SE(test_se), .CLK(CK), .Q(
        test_so36), .QN() );
  SDFFX1 DFF_594_Q_reg ( .D(g29354), .SI(test_si37), .SE(test_se), .CLK(CK), 
        .Q(g744), .QN() );
  SDFFX1 DFF_595_Q_reg ( .D(g29580), .SI(g744), .SE(test_se), .CLK(CK), .Q(
        g740), .QN() );
  SDFFX1 DFF_596_Q_reg ( .D(g13110), .SI(g740), .SE(test_se), .CLK(CK), .Q(
        g868), .QN() );
  SDFFX1 DFF_597_Q_reg ( .D(g868), .SI(g868), .SE(test_se), .CLK(CK), .Q(g5595), .QN() );
  SDFFX1 DFF_598_Q_reg ( .D(g5595), .SI(g5595), .SE(test_se), .CLK(CK), .Q(
        g869), .QN() );
  SDFFX1 DFF_599_Q_reg ( .D(n4650), .SI(g869), .SE(test_se), .CLK(CK), .Q(g963), .QN(n4363) );
  SDFFX1 DFF_600_Q_reg ( .D(g5472), .SI(g963), .SE(test_se), .CLK(CK), .Q(
        g1092), .QN(n4364) );
  SDFFX1 DFF_601_Q_reg ( .D(g6712), .SI(g1092), .SE(test_se), .CLK(CK), .Q(
        g1088), .QN(n4381) );
  SDFFX1 DFF_602_Q_reg ( .D(g5595), .SI(g1088), .SE(test_se), .CLK(CK), .Q(
        g996), .QN(n4387) );
  SDFFX1 DFF_603_Q_reg ( .D(g27257), .SI(g996), .SE(test_se), .CLK(CK), .Q(
        g1041), .QN() );
  SDFFX1 DFF_604_Q_reg ( .D(g27262), .SI(g1041), .SE(test_se), .CLK(CK), .Q(
        g1030), .QN() );
  SDFFX1 DFF_605_Q_reg ( .D(g27270), .SI(g1030), .SE(test_se), .CLK(CK), .Q(
        g1033), .QN() );
  SDFFX1 DFF_606_Q_reg ( .D(g27263), .SI(g1033), .SE(test_se), .CLK(CK), .Q(
        g1056), .QN() );
  SDFFX1 DFF_607_Q_reg ( .D(g27271), .SI(g1056), .SE(test_se), .CLK(CK), .Q(
        g1045), .QN() );
  SDFFX1 DFF_608_Q_reg ( .D(g27282), .SI(g1045), .SE(test_se), .CLK(CK), .Q(
        g1048), .QN() );
  SDFFX1 DFF_609_Q_reg ( .D(g27272), .SI(g1048), .SE(test_se), .CLK(CK), .Q(
        test_so37), .QN() );
  SDFFX1 DFF_610_Q_reg ( .D(g27283), .SI(test_si38), .SE(test_se), .CLK(CK), 
        .Q(g1060), .QN() );
  SDFFX1 DFF_611_Q_reg ( .D(g27297), .SI(g1060), .SE(test_se), .CLK(CK), .Q(
        g1063), .QN() );
  SDFFX1 DFF_612_Q_reg ( .D(g27284), .SI(g1063), .SE(test_se), .CLK(CK), .Q(
        g1085), .QN() );
  SDFFX1 DFF_613_Q_reg ( .D(g27298), .SI(g1085), .SE(test_se), .CLK(CK), .Q(
        g1075), .QN() );
  SDFFX1 DFF_614_Q_reg ( .D(g27313), .SI(g1075), .SE(test_se), .CLK(CK), .Q(
        g1078), .QN() );
  SDFFX1 DFF_615_Q_reg ( .D(g28738), .SI(g1078), .SE(test_se), .CLK(CK), .Q(
        g1095), .QN() );
  SDFFX1 DFF_616_Q_reg ( .D(g28746), .SI(g1095), .SE(test_se), .CLK(CK), .Q(
        g1098), .QN() );
  SDFFX1 DFF_617_Q_reg ( .D(g28758), .SI(g1098), .SE(test_se), .CLK(CK), .Q(
        g1101), .QN() );
  SDFFX1 DFF_618_Q_reg ( .D(g29198), .SI(g1101), .SE(test_se), .CLK(CK), .Q(
        g1104), .QN() );
  SDFFX1 DFF_619_Q_reg ( .D(g29204), .SI(g1104), .SE(test_se), .CLK(CK), .Q(
        g1107), .QN() );
  SDFFX1 DFF_620_Q_reg ( .D(g29209), .SI(g1107), .SE(test_se), .CLK(CK), .Q(
        g1110), .QN() );
  SDFFX1 DFF_621_Q_reg ( .D(g28747), .SI(g1110), .SE(test_se), .CLK(CK), .Q(
        g1114), .QN() );
  SDFFX1 DFF_622_Q_reg ( .D(g28759), .SI(g1114), .SE(test_se), .CLK(CK), .Q(
        g1115), .QN() );
  SDFFX1 DFF_623_Q_reg ( .D(g28767), .SI(g1115), .SE(test_se), .CLK(CK), .Q(
        g1113), .QN() );
  SDFFX1 DFF_624_Q_reg ( .D(g26806), .SI(g1113), .SE(test_se), .CLK(CK), .Q(
        g1116), .QN() );
  SDFFX1 DFF_625_Q_reg ( .D(g26809), .SI(g1116), .SE(test_se), .CLK(CK), .Q(
        test_so38), .QN() );
  SDFFX1 DFF_626_Q_reg ( .D(g26813), .SI(test_si39), .SE(test_se), .CLK(CK), 
        .Q(g1122), .QN() );
  SDFFX1 DFF_627_Q_reg ( .D(g26810), .SI(g1122), .SE(test_se), .CLK(CK), .Q(
        g1125), .QN() );
  SDFFX1 DFF_628_Q_reg ( .D(g26814), .SI(g1125), .SE(test_se), .CLK(CK), .Q(
        g1128), .QN() );
  SDFFX1 DFF_629_Q_reg ( .D(g26818), .SI(g1128), .SE(test_se), .CLK(CK), .Q(
        g1131), .QN() );
  SDFFX1 DFF_630_Q_reg ( .D(g27761), .SI(g1131), .SE(test_se), .CLK(CK), .Q(
        g1135), .QN() );
  SDFFX1 DFF_631_Q_reg ( .D(g27763), .SI(g1135), .SE(test_se), .CLK(CK), .Q(
        g1136), .QN() );
  SDFFX1 DFF_632_Q_reg ( .D(g27765), .SI(g1136), .SE(test_se), .CLK(CK), .Q(
        g1134), .QN() );
  SDFFX1 DFF_633_Q_reg ( .D(g29609), .SI(g1134), .SE(test_se), .CLK(CK), .Q(
        g999), .QN() );
  SDFFX1 DFF_634_Q_reg ( .D(g29612), .SI(g999), .SE(test_se), .CLK(CK), .Q(
        g1000), .QN() );
  SDFFX1 DFF_635_Q_reg ( .D(g29616), .SI(g1000), .SE(test_se), .CLK(CK), .Q(
        g1001), .QN() );
  SDFFX1 DFF_636_Q_reg ( .D(g30701), .SI(g1001), .SE(test_se), .CLK(CK), .Q(
        g1002), .QN() );
  SDFFX1 DFF_637_Q_reg ( .D(g30703), .SI(g1002), .SE(test_se), .CLK(CK), .Q(
        g1003), .QN() );
  SDFFX1 DFF_638_Q_reg ( .D(g30705), .SI(g1003), .SE(test_se), .CLK(CK), .Q(
        g1004), .QN() );
  SDFFX1 DFF_639_Q_reg ( .D(g30470), .SI(g1004), .SE(test_se), .CLK(CK), .Q(
        g1005), .QN() );
  SDFFX1 DFF_640_Q_reg ( .D(g30485), .SI(g1005), .SE(test_se), .CLK(CK), .Q(
        g1006), .QN() );
  SDFFX1 DFF_641_Q_reg ( .D(g30500), .SI(g1006), .SE(test_se), .CLK(CK), .Q(
        test_so39), .QN() );
  SDFFX1 DFF_642_Q_reg ( .D(g29170), .SI(test_si40), .SE(test_se), .CLK(CK), 
        .Q(g1009), .QN() );
  SDFFX1 DFF_643_Q_reg ( .D(g29173), .SI(g1009), .SE(test_se), .CLK(CK), .Q(
        g1010), .QN() );
  SDFFX1 DFF_644_Q_reg ( .D(g29179), .SI(g1010), .SE(test_se), .CLK(CK), .Q(
        g1008), .QN() );
  SDFFX1 DFF_645_Q_reg ( .D(g26661), .SI(g1008), .SE(test_se), .CLK(CK), .Q(
        g1090), .QN() );
  SDFFX1 DFF_646_Q_reg ( .D(g26665), .SI(g1090), .SE(test_se), .CLK(CK), .Q(
        g1091), .QN() );
  SDFFX1 DFF_647_Q_reg ( .D(g26669), .SI(g1091), .SE(test_se), .CLK(CK), .Q(
        g1089), .QN() );
  SDFFX1 DFF_648_Q_reg ( .D(n4289), .SI(g1089), .SE(test_se), .CLK(CK), .Q(
        g1137), .QN() );
  SDFFX1 DFF_649_Q_reg ( .D(g1137), .SI(g1137), .SE(test_se), .CLK(CK), .Q(
        n8027), .QN(DFF_649_n1) );
  SDFFX1 DFF_650_Q_reg ( .D(n4567), .SI(n8027), .SE(test_se), .CLK(CK), .Q(
        g1139), .QN() );
  SDFFX1 DFF_651_Q_reg ( .D(g1139), .SI(g1139), .SE(test_se), .CLK(CK), .Q(
        n8026), .QN(DFF_651_n1) );
  SDFFX1 DFF_652_Q_reg ( .D(n4559), .SI(n8026), .SE(test_se), .CLK(CK), .Q(
        g1141), .QN() );
  SDFFX1 DFF_653_Q_reg ( .D(g1141), .SI(g1141), .SE(test_se), .CLK(CK), .Q(
        n8025), .QN(DFF_653_n1) );
  SDFFX1 DFF_654_Q_reg ( .D(n4327), .SI(n8025), .SE(test_se), .CLK(CK), .Q(
        g967), .QN() );
  SDFFX1 DFF_655_Q_reg ( .D(g967), .SI(g967), .SE(test_se), .CLK(CK), .Q(n8024), .QN(DFF_655_n1) );
  SDFFX1 DFF_656_Q_reg ( .D(n4391), .SI(n8024), .SE(test_se), .CLK(CK), .Q(
        g969), .QN() );
  SDFFX1 DFF_657_Q_reg ( .D(g969), .SI(g969), .SE(test_se), .CLK(CK), .Q(
        test_so40), .QN(DFF_657_n1) );
  SDFFX1 DFF_658_Q_reg ( .D(n4321), .SI(test_si41), .SE(test_se), .CLK(CK), 
        .Q(g971), .QN() );
  SDFFX1 DFF_659_Q_reg ( .D(g971), .SI(g971), .SE(test_se), .CLK(CK), .Q(n8021), .QN(DFF_659_n1) );
  SDFFX1 DFF_660_Q_reg ( .D(n4375), .SI(n8021), .SE(test_se), .CLK(CK), .Q(
        g973), .QN() );
  SDFFX1 DFF_661_Q_reg ( .D(g973), .SI(g973), .SE(test_se), .CLK(CK), .Q(n8020), .QN(DFF_661_n1) );
  SDFFX1 DFF_662_Q_reg ( .D(n4379), .SI(n8020), .SE(test_se), .CLK(CK), .Q(
        g975), .QN() );
  SDFFX1 DFF_663_Q_reg ( .D(g975), .SI(g975), .SE(test_se), .CLK(CK), .Q(n8019), .QN(DFF_663_n1) );
  SDFFX1 DFF_664_Q_reg ( .D(g2873), .SI(n8019), .SE(test_se), .CLK(CK), .Q(
        g977), .QN() );
  SDFFX1 DFF_665_Q_reg ( .D(g977), .SI(g977), .SE(test_se), .CLK(CK), .Q(n8018), .QN(n4486) );
  SDFFX1 DFF_666_Q_reg ( .D(n4283), .SI(n8018), .SE(test_se), .CLK(CK), .Q(
        g986), .QN(n4432) );
  SDFFX1 DFF_667_Q_reg ( .D(g26183), .SI(g986), .SE(test_se), .CLK(CK), .Q(
        g992), .QN() );
  SDFFX1 DFF_678_Q_reg ( .D(n4277), .SI(g992), .SE(test_se), .CLK(CK), .Q(
        n8017), .QN(n4583) );
  SDFFX1 DFF_679_Q_reg ( .D(g1041), .SI(n8017), .SE(test_se), .CLK(CK), .Q(
        g1029), .QN() );
  SDFFX1 DFF_680_Q_reg ( .D(g1029), .SI(g1029), .SE(test_se), .CLK(CK), .Q(
        g1036), .QN() );
  SDFFX1 DFF_681_Q_reg ( .D(g1030), .SI(g1036), .SE(test_se), .CLK(CK), .Q(
        g1037), .QN() );
  SDFFX1 DFF_682_Q_reg ( .D(g1037), .SI(g1037), .SE(test_se), .CLK(CK), .Q(
        g1038), .QN() );
  SDFFX1 DFF_683_Q_reg ( .D(g1033), .SI(g1038), .SE(test_se), .CLK(CK), .Q(
        test_so41), .QN() );
  SDFFX1 DFF_684_Q_reg ( .D(test_so41), .SI(test_si42), .SE(test_se), .CLK(CK), 
        .Q(g1040), .QN() );
  SDFFX1 DFF_685_Q_reg ( .D(g1056), .SI(g1040), .SE(test_se), .CLK(CK), .Q(
        g1044), .QN() );
  SDFFX1 DFF_686_Q_reg ( .D(g1044), .SI(g1044), .SE(test_se), .CLK(CK), .Q(
        g1051), .QN() );
  SDFFX1 DFF_687_Q_reg ( .D(g1045), .SI(g1051), .SE(test_se), .CLK(CK), .Q(
        g1052), .QN() );
  SDFFX1 DFF_688_Q_reg ( .D(g1052), .SI(g1052), .SE(test_se), .CLK(CK), .Q(
        g1053), .QN() );
  SDFFX1 DFF_689_Q_reg ( .D(g1048), .SI(g1053), .SE(test_se), .CLK(CK), .Q(
        g1054), .QN() );
  SDFFX1 DFF_690_Q_reg ( .D(g1054), .SI(g1054), .SE(test_se), .CLK(CK), .Q(
        g1055), .QN() );
  SDFFX1 DFF_691_Q_reg ( .D(test_so37), .SI(g1055), .SE(test_se), .CLK(CK), 
        .Q(g1059), .QN() );
  SDFFX1 DFF_692_Q_reg ( .D(g1059), .SI(g1059), .SE(test_se), .CLK(CK), .Q(
        g1066), .QN() );
  SDFFX1 DFF_693_Q_reg ( .D(g1060), .SI(g1066), .SE(test_se), .CLK(CK), .Q(
        g1067), .QN() );
  SDFFX1 DFF_694_Q_reg ( .D(g1067), .SI(g1067), .SE(test_se), .CLK(CK), .Q(
        g1068), .QN() );
  SDFFX1 DFF_695_Q_reg ( .D(g1063), .SI(g1068), .SE(test_se), .CLK(CK), .Q(
        g1069), .QN() );
  SDFFX1 DFF_696_Q_reg ( .D(g1069), .SI(g1069), .SE(test_se), .CLK(CK), .Q(
        g1070), .QN() );
  SDFFX1 DFF_697_Q_reg ( .D(g1085), .SI(g1070), .SE(test_se), .CLK(CK), .Q(
        g1074), .QN() );
  SDFFX1 DFF_698_Q_reg ( .D(g1074), .SI(g1074), .SE(test_se), .CLK(CK), .Q(
        g1081), .QN() );
  SDFFX1 DFF_699_Q_reg ( .D(g1075), .SI(g1081), .SE(test_se), .CLK(CK), .Q(
        test_so42), .QN() );
  SDFFX1 DFF_700_Q_reg ( .D(test_so42), .SI(test_si43), .SE(test_se), .CLK(CK), 
        .Q(g1083), .QN() );
  SDFFX1 DFF_701_Q_reg ( .D(g1078), .SI(g1083), .SE(test_se), .CLK(CK), .Q(
        g1084), .QN() );
  SDFFX1 DFF_702_Q_reg ( .D(g1084), .SI(g1084), .SE(test_se), .CLK(CK), .Q(
        g1011), .QN() );
  SDFFX1 DFF_703_Q_reg ( .D(n4598), .SI(g1011), .SE(test_se), .CLK(CK), .Q(
        g5657), .QN() );
  SDFFX1 DFF_704_Q_reg ( .D(g5657), .SI(g5657), .SE(test_se), .CLK(CK), .Q(
        g5686), .QN() );
  SDFFX1 DFF_705_Q_reg ( .D(g5686), .SI(g5686), .SE(test_se), .CLK(CK), .Q(
        g1024), .QN() );
  SDFFX1 DFF_706_Q_reg ( .D(n4598), .SI(g1024), .SE(test_se), .CLK(CK), .Q(
        g1231), .QN(n4371) );
  SDFFX1 DFF_707_Q_reg ( .D(g6750), .SI(g1231), .SE(test_se), .CLK(CK), .Q(
        g1237), .QN(n4316) );
  SDFFX1 DFF_708_Q_reg ( .D(n4626), .SI(g1237), .SE(test_se), .CLK(CK), .Q(
        g1236), .QN(n4300) );
  SDFFX1 DFF_709_Q_reg ( .D(g21843), .SI(g1236), .SE(test_se), .CLK(CK), .Q(
        g1240), .QN() );
  SDFFX1 DFF_710_Q_reg ( .D(g18707), .SI(g1240), .SE(test_se), .CLK(CK), .Q(
        g1243), .QN(n4353) );
  SDFFX1 DFF_711_Q_reg ( .D(g18763), .SI(g1243), .SE(test_se), .CLK(CK), .Q(
        g1196), .QN(n4304) );
  SDFFX1 DFF_712_Q_reg ( .D(g12507), .SI(g1196), .SE(test_se), .CLK(CK), .Q(
        g1199), .QN() );
  SDFFX1 DFF_713_Q_reg ( .D(g1199), .SI(g1199), .SE(test_se), .CLK(CK), .Q(
        g1209), .QN() );
  SDFFX1 DFF_714_Q_reg ( .D(g1209), .SI(g1209), .SE(test_se), .CLK(CK), .Q(
        g1210), .QN() );
  SDFFX1 DFF_715_Q_reg ( .D(g1142), .SI(g1210), .SE(test_se), .CLK(CK), .Q(
        test_so43), .QN() );
  SDFFX1 DFF_716_Q_reg ( .D(test_so43), .SI(test_si44), .SE(test_se), .CLK(CK), 
        .Q(g1255), .QN() );
  SDFFX1 DFF_717_Q_reg ( .D(g1145), .SI(g1255), .SE(test_se), .CLK(CK), .Q(
        g1256), .QN() );
  SDFFX1 DFF_718_Q_reg ( .D(g1256), .SI(g1256), .SE(test_se), .CLK(CK), .Q(
        g1257), .QN() );
  SDFFX1 DFF_719_Q_reg ( .D(g1148), .SI(g1257), .SE(test_se), .CLK(CK), .Q(
        g1258), .QN() );
  SDFFX1 DFF_720_Q_reg ( .D(g1258), .SI(g1258), .SE(test_se), .CLK(CK), .Q(
        g1259), .QN() );
  SDFFX1 DFF_721_Q_reg ( .D(g1152), .SI(g1259), .SE(test_se), .CLK(CK), .Q(
        g1260), .QN() );
  SDFFX1 DFF_722_Q_reg ( .D(g1260), .SI(g1260), .SE(test_se), .CLK(CK), .Q(
        g1251), .QN() );
  SDFFX1 DFF_723_Q_reg ( .D(g1155), .SI(g1251), .SE(test_se), .CLK(CK), .Q(
        g1252), .QN() );
  SDFFX1 DFF_724_Q_reg ( .D(g1252), .SI(g1252), .SE(test_se), .CLK(CK), .Q(
        g1253), .QN() );
  SDFFX1 DFF_725_Q_reg ( .D(g1158), .SI(g1253), .SE(test_se), .CLK(CK), .Q(
        g1254), .QN() );
  SDFFX1 DFF_726_Q_reg ( .D(g1254), .SI(g1254), .SE(test_se), .CLK(CK), .Q(
        g1176), .QN() );
  SDFFX1 DFF_727_Q_reg ( .D(n4650), .SI(g1176), .SE(test_se), .CLK(CK), .Q(
        g7961), .QN(n4460) );
  SDFFX1 DFF_728_Q_reg ( .D(g7961), .SI(g7961), .SE(test_se), .CLK(CK), .Q(
        g8007), .QN(n4459) );
  SDFFX1 DFF_729_Q_reg ( .D(g8007), .SI(g8007), .SE(test_se), .CLK(CK), .Q(
        g1172), .QN(n4465) );
  SDFFX1 DFF_730_Q_reg ( .D(g23081), .SI(g1172), .SE(test_se), .CLK(CK), .Q(
        g1173), .QN() );
  SDFFX1 DFF_731_Q_reg ( .D(g23111), .SI(g1173), .SE(test_se), .CLK(CK), .Q(
        test_so44), .QN() );
  SDFFX1 DFF_732_Q_reg ( .D(g23126), .SI(test_si45), .SE(test_se), .CLK(CK), 
        .Q(g1175), .QN() );
  SDFFX1 DFF_733_Q_reg ( .D(g23392), .SI(g1175), .SE(test_se), .CLK(CK), .Q(
        g1142), .QN() );
  SDFFX1 DFF_734_Q_reg ( .D(g23406), .SI(g1142), .SE(test_se), .CLK(CK), .Q(
        g1145), .QN() );
  SDFFX1 DFF_735_Q_reg ( .D(g24179), .SI(g1145), .SE(test_se), .CLK(CK), .Q(
        g1148), .QN() );
  SDFFX1 DFF_736_Q_reg ( .D(g24181), .SI(g1148), .SE(test_se), .CLK(CK), .Q(
        g1164), .QN() );
  SDFFX1 DFF_737_Q_reg ( .D(g24213), .SI(g1164), .SE(test_se), .CLK(CK), .Q(
        g1165), .QN() );
  SDFFX1 DFF_738_Q_reg ( .D(g24223), .SI(g1165), .SE(test_se), .CLK(CK), .Q(
        g1166), .QN() );
  SDFFX1 DFF_739_Q_reg ( .D(g23110), .SI(g1166), .SE(test_se), .CLK(CK), .Q(
        g1167), .QN() );
  SDFFX1 DFF_740_Q_reg ( .D(g23014), .SI(g1167), .SE(test_se), .CLK(CK), .Q(
        g1171), .QN() );
  SDFFX1 DFF_741_Q_reg ( .D(g23039), .SI(g1171), .SE(test_se), .CLK(CK), .Q(
        g1151), .QN() );
  SDFFX1 DFF_742_Q_reg ( .D(g24212), .SI(g1151), .SE(test_se), .CLK(CK), .Q(
        g1152), .QN() );
  SDFFX1 DFF_743_Q_reg ( .D(g24222), .SI(g1152), .SE(test_se), .CLK(CK), .Q(
        g1155), .QN() );
  SDFFX1 DFF_744_Q_reg ( .D(g24235), .SI(g1155), .SE(test_se), .CLK(CK), .Q(
        g1158), .QN() );
  SDFFX1 DFF_745_Q_reg ( .D(g12467), .SI(g1158), .SE(test_se), .CLK(CK), .Q(
        g1214), .QN() );
  SDFFX1 DFF_746_Q_reg ( .D(g1214), .SI(g1214), .SE(test_se), .CLK(CK), .Q(
        g1221), .QN() );
  SDFFX1 DFF_747_Q_reg ( .D(g1221), .SI(g1221), .SE(test_se), .CLK(CK), .Q(
        test_so45), .QN() );
  SDFFX1 DFF_748_Q_reg ( .D(g13155), .SI(test_si46), .SE(test_se), .CLK(CK), 
        .Q(g1229), .QN() );
  SDFFX1 DFF_749_Q_reg ( .D(g1229), .SI(g1229), .SE(test_se), .CLK(CK), .Q(
        n4549), .QN() );
  SDFFX1 DFF_750_Q_reg ( .D(n1817), .SI(n4549), .SE(test_se), .CLK(CK), .Q(
        n4361), .QN() );
  SDFFX1 DFF_751_Q_reg ( .D(g13124), .SI(n4361), .SE(test_se), .CLK(CK), .Q(
        g1235), .QN() );
  SDFFX1 DFF_752_Q_reg ( .D(g1235), .SI(g1235), .SE(test_se), .CLK(CK), .Q(
        g1186), .QN(n4548) );
  SDFFX1 DFF_753_Q_reg ( .D(g13171), .SI(g1186), .SE(test_se), .CLK(CK), .Q(
        g1244), .QN() );
  SDFFX1 DFF_754_Q_reg ( .D(g1244), .SI(g1244), .SE(test_se), .CLK(CK), .Q(
        g1245), .QN() );
  SDFFX1 DFF_755_Q_reg ( .D(g27273), .SI(g1245), .SE(test_se), .CLK(CK), .Q(
        g1262), .QN() );
  SDFFX1 DFF_756_Q_reg ( .D(g27285), .SI(g1262), .SE(test_se), .CLK(CK), .Q(
        g1263), .QN() );
  SDFFX1 DFF_757_Q_reg ( .D(g27299), .SI(g1263), .SE(test_se), .CLK(CK), .Q(
        g1261), .QN() );
  SDFFX1 DFF_758_Q_reg ( .D(g27286), .SI(g1261), .SE(test_se), .CLK(CK), .Q(
        g1265), .QN() );
  SDFFX1 DFF_759_Q_reg ( .D(g27300), .SI(g1265), .SE(test_se), .CLK(CK), .Q(
        g1266), .QN() );
  SDFFX1 DFF_760_Q_reg ( .D(g27314), .SI(g1266), .SE(test_se), .CLK(CK), .Q(
        g1264), .QN() );
  SDFFX1 DFF_761_Q_reg ( .D(g27301), .SI(g1264), .SE(test_se), .CLK(CK), .Q(
        g1268), .QN() );
  SDFFX1 DFF_762_Q_reg ( .D(g27315), .SI(g1268), .SE(test_se), .CLK(CK), .Q(
        g1269), .QN() );
  SDFFX1 DFF_763_Q_reg ( .D(g27328), .SI(g1269), .SE(test_se), .CLK(CK), .Q(
        test_so46), .QN() );
  SDFFX1 DFF_764_Q_reg ( .D(g27316), .SI(test_si47), .SE(test_se), .CLK(CK), 
        .Q(g1271), .QN() );
  SDFFX1 DFF_765_Q_reg ( .D(g27329), .SI(g1271), .SE(test_se), .CLK(CK), .Q(
        g1272), .QN() );
  SDFFX1 DFF_766_Q_reg ( .D(g27339), .SI(g1272), .SE(test_se), .CLK(CK), .Q(
        g1270), .QN() );
  SDFFX1 DFF_767_Q_reg ( .D(g24501), .SI(g1270), .SE(test_se), .CLK(CK), .Q(
        g1273), .QN() );
  SDFFX1 DFF_768_Q_reg ( .D(g24510), .SI(g1273), .SE(test_se), .CLK(CK), .Q(
        g1276), .QN() );
  SDFFX1 DFF_769_Q_reg ( .D(g24521), .SI(g1276), .SE(test_se), .CLK(CK), .Q(
        g1279), .QN() );
  SDFFX1 DFF_770_Q_reg ( .D(g24511), .SI(g1279), .SE(test_se), .CLK(CK), .Q(
        g1282), .QN() );
  SDFFX1 DFF_771_Q_reg ( .D(g24522), .SI(g1282), .SE(test_se), .CLK(CK), .Q(
        g1285), .QN() );
  SDFFX1 DFF_772_Q_reg ( .D(g24532), .SI(g1285), .SE(test_se), .CLK(CK), .Q(
        g1288), .QN() );
  SDFFX1 DFF_773_Q_reg ( .D(g28351), .SI(g1288), .SE(test_se), .CLK(CK), .Q(
        g1300), .QN() );
  SDFFX1 DFF_774_Q_reg ( .D(g28355), .SI(g1300), .SE(test_se), .CLK(CK), .Q(
        g1303), .QN() );
  SDFFX1 DFF_775_Q_reg ( .D(g28360), .SI(g1303), .SE(test_se), .CLK(CK), .Q(
        g1306), .QN() );
  SDFFX1 DFF_776_Q_reg ( .D(g28346), .SI(g1306), .SE(test_se), .CLK(CK), .Q(
        g1291), .QN() );
  SDFFX1 DFF_777_Q_reg ( .D(g28350), .SI(g1291), .SE(test_se), .CLK(CK), .Q(
        g1294), .QN() );
  SDFFX1 DFF_778_Q_reg ( .D(g28354), .SI(g1294), .SE(test_se), .CLK(CK), .Q(
        g1297), .QN() );
  SDFFX1 DFF_779_Q_reg ( .D(g26547), .SI(g1297), .SE(test_se), .CLK(CK), .Q(
        test_so47), .QN() );
  SDFFX1 DFF_780_Q_reg ( .D(g26557), .SI(test_si48), .SE(test_se), .CLK(CK), 
        .Q(g1180), .QN() );
  SDFFX1 DFF_781_Q_reg ( .D(g26569), .SI(g1180), .SE(test_se), .CLK(CK), .Q(
        g1183), .QN() );
  SDFFX1 DFF_782_Q_reg ( .D(g1186), .SI(g1183), .SE(test_se), .CLK(CK), .Q(
        g1192), .QN(n4454) );
  SDFFX1 DFF_783_Q_reg ( .D(g22615), .SI(g1192), .SE(test_se), .CLK(CK), .Q(
        n8009), .QN(DFF_783_n1) );
  SDFFX1 DFF_792_Q_reg ( .D(n1829), .SI(n8009), .SE(test_se), .CLK(CK), .Q(
        g16355), .QN(DFF_792_n1) );
  SDFFX1 DFF_793_Q_reg ( .D(g16355), .SI(g16355), .SE(test_se), .CLK(CK), .Q(
        g1211), .QN() );
  SDFFX1 DFF_794_Q_reg ( .D(DFF_649_n1), .SI(g1211), .SE(test_se), .CLK(CK), 
        .Q(n8008), .QN(DFF_794_n1) );
  SDFFX1 DFF_795_Q_reg ( .D(DFF_651_n1), .SI(n8008), .SE(test_se), .CLK(CK), 
        .Q(n8007), .QN(DFF_795_n1) );
  SDFFX1 DFF_796_Q_reg ( .D(DFF_653_n1), .SI(n8007), .SE(test_se), .CLK(CK), 
        .Q(n8006), .QN(DFF_796_n1) );
  SDFFX1 DFF_797_Q_reg ( .D(DFF_655_n1), .SI(n8006), .SE(test_se), .CLK(CK), 
        .Q(n8005), .QN(DFF_797_n1) );
  SDFFX1 DFF_798_Q_reg ( .D(DFF_657_n1), .SI(n8005), .SE(test_se), .CLK(CK), 
        .Q(n8004), .QN(DFF_798_n1) );
  SDFFX1 DFF_799_Q_reg ( .D(DFF_659_n1), .SI(n8004), .SE(test_se), .CLK(CK), 
        .Q(n8003), .QN(DFF_799_n1) );
  SDFFX1 DFF_800_Q_reg ( .D(DFF_661_n1), .SI(n8003), .SE(test_se), .CLK(CK), 
        .Q(g1222), .QN() );
  SDFFX1 DFF_801_Q_reg ( .D(DFF_663_n1), .SI(g1222), .SE(test_se), .CLK(CK), 
        .Q(g1223), .QN() );
  SDFFX1 DFF_802_Q_reg ( .D(g24072), .SI(g1223), .SE(test_se), .CLK(CK), .Q(
        g1224), .QN(n4489) );
  SDFFX1 DFF_803_Q_reg ( .D(n4486), .SI(g1224), .SE(test_se), .CLK(CK), .Q(
        test_so48), .QN(DFF_803_n1) );
  SDFFX1 DFF_805_Q_reg ( .D(g6979), .SI(g6979), .SE(test_se), .CLK(CK), .Q(
        g7161), .QN(n4358) );
  SDFFX1 DFF_806_Q_reg ( .D(g7161), .SI(g7161), .SE(test_se), .CLK(CK), .Q(
        g1315), .QN(n4294) );
  SDFFX1 DFF_807_Q_reg ( .D(g16671), .SI(g1315), .SE(test_se), .CLK(CK), .Q(
        g1316), .QN() );
  SDFFX1 DFF_808_Q_reg ( .D(g20333), .SI(g1316), .SE(test_se), .CLK(CK), .Q(
        g1345), .QN(n4428) );
  SDFFX1 DFF_809_Q_reg ( .D(g20717), .SI(g1345), .SE(test_se), .CLK(CK), .Q(
        g1326), .QN(n4402) );
  SDFFX1 DFF_810_Q_reg ( .D(g21969), .SI(g1326), .SE(test_se), .CLK(CK), .Q(
        g1319), .QN(n4476) );
  SDFFX1 DFF_811_Q_reg ( .D(g23329), .SI(g1319), .SE(test_se), .CLK(CK), .Q(
        g1339), .QN(n4421) );
  SDFFX1 DFF_812_Q_reg ( .D(g24430), .SI(g1339), .SE(test_se), .CLK(CK), .Q(
        g1332), .QN(n4412) );
  SDFFX1 DFF_813_Q_reg ( .D(g25189), .SI(g1332), .SE(test_se), .CLK(CK), .Q(
        g1346), .QN(n4401) );
  SDFFX1 DFF_814_Q_reg ( .D(g26666), .SI(g1346), .SE(test_se), .CLK(CK), .Q(
        g1358), .QN(n4411) );
  SDFFX1 DFF_815_Q_reg ( .D(g26781), .SI(g1358), .SE(test_se), .CLK(CK), .Q(
        g1352), .QN(n4469) );
  SDFFX1 DFF_816_Q_reg ( .D(g27678), .SI(g1352), .SE(test_se), .CLK(CK), .Q(
        g1365), .QN(n4475) );
  SDFFX1 DFF_817_Q_reg ( .D(g27718), .SI(g1365), .SE(test_se), .CLK(CK), .Q(
        g1372), .QN(n4395) );
  SDFFX1 DFF_818_Q_reg ( .D(g28321), .SI(g1372), .SE(test_se), .CLK(CK), .Q(
        g1378), .QN(n4417) );
  SDFFX1 DFF_819_Q_reg ( .D(g20882), .SI(g1378), .SE(test_se), .CLK(CK), .Q(
        test_so49), .QN() );
  SDFFX1 DFF_820_Q_reg ( .D(g20896), .SI(test_si50), .SE(test_se), .CLK(CK), 
        .Q(g1386), .QN() );
  SDFFX1 DFF_821_Q_reg ( .D(g20910), .SI(g1386), .SE(test_se), .CLK(CK), .Q(
        g1384), .QN() );
  SDFFX1 DFF_822_Q_reg ( .D(g20897), .SI(g1384), .SE(test_se), .CLK(CK), .Q(
        g1388), .QN() );
  SDFFX1 DFF_823_Q_reg ( .D(g20911), .SI(g1388), .SE(test_se), .CLK(CK), .Q(
        g1389), .QN() );
  SDFFX1 DFF_824_Q_reg ( .D(g20925), .SI(g1389), .SE(test_se), .CLK(CK), .Q(
        g1387), .QN() );
  SDFFX1 DFF_825_Q_reg ( .D(g20912), .SI(g1387), .SE(test_se), .CLK(CK), .Q(
        g1391), .QN() );
  SDFFX1 DFF_826_Q_reg ( .D(g20926), .SI(g1391), .SE(test_se), .CLK(CK), .Q(
        g1392), .QN() );
  SDFFX1 DFF_827_Q_reg ( .D(g20949), .SI(g1392), .SE(test_se), .CLK(CK), .Q(
        g1390), .QN() );
  SDFFX1 DFF_828_Q_reg ( .D(g20927), .SI(g1390), .SE(test_se), .CLK(CK), .Q(
        g1394), .QN() );
  SDFFX1 DFF_829_Q_reg ( .D(g20950), .SI(g1394), .SE(test_se), .CLK(CK), .Q(
        g1395), .QN() );
  SDFFX1 DFF_830_Q_reg ( .D(g20972), .SI(g1395), .SE(test_se), .CLK(CK), .Q(
        g1393), .QN() );
  SDFFX1 DFF_831_Q_reg ( .D(g20951), .SI(g1393), .SE(test_se), .CLK(CK), .Q(
        g1397), .QN() );
  SDFFX1 DFF_832_Q_reg ( .D(g20973), .SI(g1397), .SE(test_se), .CLK(CK), .Q(
        g1398), .QN() );
  SDFFX1 DFF_833_Q_reg ( .D(g20993), .SI(g1398), .SE(test_se), .CLK(CK), .Q(
        g1396), .QN() );
  SDFFX1 DFF_834_Q_reg ( .D(g20974), .SI(g1396), .SE(test_se), .CLK(CK), .Q(
        g1400), .QN() );
  SDFFX1 DFF_835_Q_reg ( .D(g20994), .SI(g1400), .SE(test_se), .CLK(CK), .Q(
        test_so50), .QN() );
  SDFFX1 DFF_836_Q_reg ( .D(g21015), .SI(test_si51), .SE(test_se), .CLK(CK), 
        .Q(g1399), .QN() );
  SDFFX1 DFF_837_Q_reg ( .D(g20995), .SI(g1399), .SE(test_se), .CLK(CK), .Q(
        g1403), .QN() );
  SDFFX1 DFF_838_Q_reg ( .D(g21016), .SI(g1403), .SE(test_se), .CLK(CK), .Q(
        g1404), .QN() );
  SDFFX1 DFF_839_Q_reg ( .D(g21033), .SI(g1404), .SE(test_se), .CLK(CK), .Q(
        g1402), .QN() );
  SDFFX1 DFF_840_Q_reg ( .D(g21017), .SI(g1402), .SE(test_se), .CLK(CK), .Q(
        g1406), .QN() );
  SDFFX1 DFF_841_Q_reg ( .D(g21034), .SI(g1406), .SE(test_se), .CLK(CK), .Q(
        g1407), .QN() );
  SDFFX1 DFF_842_Q_reg ( .D(g21052), .SI(g1407), .SE(test_se), .CLK(CK), .Q(
        g1405), .QN() );
  SDFFX1 DFF_843_Q_reg ( .D(g21035), .SI(g1405), .SE(test_se), .CLK(CK), .Q(
        g1409), .QN() );
  SDFFX1 DFF_844_Q_reg ( .D(g21053), .SI(g1409), .SE(test_se), .CLK(CK), .Q(
        g1410), .QN() );
  SDFFX1 DFF_845_Q_reg ( .D(g21070), .SI(g1410), .SE(test_se), .CLK(CK), .Q(
        g1408), .QN() );
  SDFFX1 DFF_846_Q_reg ( .D(g20883), .SI(g1408), .SE(test_se), .CLK(CK), .Q(
        g1412), .QN() );
  SDFFX1 DFF_847_Q_reg ( .D(g20898), .SI(g1412), .SE(test_se), .CLK(CK), .Q(
        g1413), .QN() );
  SDFFX1 DFF_848_Q_reg ( .D(g20913), .SI(g1413), .SE(test_se), .CLK(CK), .Q(
        g1411), .QN() );
  SDFFX1 DFF_849_Q_reg ( .D(g20952), .SI(g1411), .SE(test_se), .CLK(CK), .Q(
        g1415), .QN() );
  SDFFX1 DFF_850_Q_reg ( .D(g20975), .SI(g1415), .SE(test_se), .CLK(CK), .Q(
        g1416), .QN() );
  SDFFX1 DFF_851_Q_reg ( .D(g20996), .SI(g1416), .SE(test_se), .CLK(CK), .Q(
        test_so51), .QN() );
  SDFFX1 DFF_852_Q_reg ( .D(g20976), .SI(test_si52), .SE(test_se), .CLK(CK), 
        .Q(g1418), .QN() );
  SDFFX1 DFF_853_Q_reg ( .D(g20997), .SI(g1418), .SE(test_se), .CLK(CK), .Q(
        g1419), .QN() );
  SDFFX1 DFF_854_Q_reg ( .D(g21018), .SI(g1419), .SE(test_se), .CLK(CK), .Q(
        g1417), .QN() );
  SDFFX1 DFF_855_Q_reg ( .D(g25263), .SI(g1417), .SE(test_se), .CLK(CK), .Q(
        g1421), .QN() );
  SDFFX1 DFF_856_Q_reg ( .D(g25267), .SI(g1421), .SE(test_se), .CLK(CK), .Q(
        g1422), .QN() );
  SDFFX1 DFF_857_Q_reg ( .D(g25270), .SI(g1422), .SE(test_se), .CLK(CK), .Q(
        g1420), .QN() );
  SDFFX1 DFF_858_Q_reg ( .D(g22234), .SI(g1420), .SE(test_se), .CLK(CK), .Q(
        g1424), .QN() );
  SDFFX1 DFF_859_Q_reg ( .D(g22247), .SI(g1424), .SE(test_se), .CLK(CK), .Q(
        g1425), .QN() );
  SDFFX1 DFF_860_Q_reg ( .D(g22263), .SI(g1425), .SE(test_se), .CLK(CK), .Q(
        g1423), .QN() );
  SDFFX1 DFF_861_Q_reg ( .D(n4650), .SI(g1423), .SE(test_se), .CLK(CK), .Q(
        g1520), .QN(n4317) );
  SDFFX1 DFF_862_Q_reg ( .D(g6573), .SI(g1520), .SE(test_se), .CLK(CK), .Q(
        g6782), .QN(n4515) );
  SDFFX1 DFF_863_Q_reg ( .D(n4589), .SI(g6782), .SE(test_se), .CLK(CK), .Q(
        g1547), .QN(n4368) );
  SDFFX1 DFF_864_Q_reg ( .D(g22149), .SI(g1547), .SE(test_se), .CLK(CK), .Q(
        g1512), .QN() );
  SDFFX1 DFF_865_Q_reg ( .D(g22166), .SI(g1512), .SE(test_se), .CLK(CK), .Q(
        g1513), .QN() );
  SDFFX1 DFF_866_Q_reg ( .D(g22178), .SI(g1513), .SE(test_se), .CLK(CK), .Q(
        g1511), .QN() );
  SDFFX1 DFF_867_Q_reg ( .D(g22167), .SI(g1511), .SE(test_se), .CLK(CK), .Q(
        test_so52), .QN() );
  SDFFX1 DFF_868_Q_reg ( .D(g22179), .SI(test_si53), .SE(test_se), .CLK(CK), 
        .Q(g1516), .QN() );
  SDFFX1 DFF_869_Q_reg ( .D(g22191), .SI(g1516), .SE(test_se), .CLK(CK), .Q(
        g1514), .QN() );
  SDFFX1 DFF_870_Q_reg ( .D(g22035), .SI(g1514), .SE(test_se), .CLK(CK), .Q(
        g1524), .QN() );
  SDFFX1 DFF_871_Q_reg ( .D(g22043), .SI(g1524), .SE(test_se), .CLK(CK), .Q(
        g1525), .QN() );
  SDFFX1 DFF_872_Q_reg ( .D(g22057), .SI(g1525), .SE(test_se), .CLK(CK), .Q(
        g1523), .QN() );
  SDFFX1 DFF_873_Q_reg ( .D(g22044), .SI(g1523), .SE(test_se), .CLK(CK), .Q(
        g1527), .QN() );
  SDFFX1 DFF_874_Q_reg ( .D(g22058), .SI(g1527), .SE(test_se), .CLK(CK), .Q(
        g1528), .QN() );
  SDFFX1 DFF_875_Q_reg ( .D(g22073), .SI(g1528), .SE(test_se), .CLK(CK), .Q(
        g1526), .QN() );
  SDFFX1 DFF_876_Q_reg ( .D(g22059), .SI(g1526), .SE(test_se), .CLK(CK), .Q(
        g1530), .QN() );
  SDFFX1 DFF_877_Q_reg ( .D(g22074), .SI(g1530), .SE(test_se), .CLK(CK), .Q(
        g1531), .QN() );
  SDFFX1 DFF_878_Q_reg ( .D(g22090), .SI(g1531), .SE(test_se), .CLK(CK), .Q(
        g1529), .QN() );
  SDFFX1 DFF_879_Q_reg ( .D(g22075), .SI(g1529), .SE(test_se), .CLK(CK), .Q(
        g1533), .QN() );
  SDFFX1 DFF_880_Q_reg ( .D(g22091), .SI(g1533), .SE(test_se), .CLK(CK), .Q(
        g1534), .QN() );
  SDFFX1 DFF_881_Q_reg ( .D(g22112), .SI(g1534), .SE(test_se), .CLK(CK), .Q(
        g1532), .QN() );
  SDFFX1 DFF_882_Q_reg ( .D(g22092), .SI(g1532), .SE(test_se), .CLK(CK), .Q(
        g1536), .QN() );
  SDFFX1 DFF_883_Q_reg ( .D(g22113), .SI(g1536), .SE(test_se), .CLK(CK), .Q(
        test_so53), .QN() );
  SDFFX1 DFF_884_Q_reg ( .D(g22130), .SI(test_si54), .SE(test_se), .CLK(CK), 
        .Q(g1535), .QN() );
  SDFFX1 DFF_885_Q_reg ( .D(g22114), .SI(g1535), .SE(test_se), .CLK(CK), .Q(
        g1539), .QN() );
  SDFFX1 DFF_886_Q_reg ( .D(g22131), .SI(g1539), .SE(test_se), .CLK(CK), .Q(
        g1540), .QN() );
  SDFFX1 DFF_887_Q_reg ( .D(g22150), .SI(g1540), .SE(test_se), .CLK(CK), .Q(
        g1538), .QN() );
  SDFFX1 DFF_888_Q_reg ( .D(g22132), .SI(g1538), .SE(test_se), .CLK(CK), .Q(
        g1542), .QN() );
  SDFFX1 DFF_889_Q_reg ( .D(g22151), .SI(g1542), .SE(test_se), .CLK(CK), .Q(
        g1543), .QN() );
  SDFFX1 DFF_890_Q_reg ( .D(g22168), .SI(g1543), .SE(test_se), .CLK(CK), .Q(
        g1541), .QN() );
  SDFFX1 DFF_891_Q_reg ( .D(g22152), .SI(g1541), .SE(test_se), .CLK(CK), .Q(
        g1545), .QN() );
  SDFFX1 DFF_892_Q_reg ( .D(g22169), .SI(g1545), .SE(test_se), .CLK(CK), .Q(
        g1546), .QN() );
  SDFFX1 DFF_893_Q_reg ( .D(g22180), .SI(g1546), .SE(test_se), .CLK(CK), .Q(
        g1544), .QN() );
  SDFFX1 DFF_894_Q_reg ( .D(g25217), .SI(g1544), .SE(test_se), .CLK(CK), .Q(
        g1551), .QN() );
  SDFFX1 DFF_895_Q_reg ( .D(g25224), .SI(g1551), .SE(test_se), .CLK(CK), .Q(
        g1552), .QN() );
  SDFFX1 DFF_896_Q_reg ( .D(g25233), .SI(g1552), .SE(test_se), .CLK(CK), .Q(
        g1550), .QN() );
  SDFFX1 DFF_897_Q_reg ( .D(g25225), .SI(g1550), .SE(test_se), .CLK(CK), .Q(
        g1554), .QN() );
  SDFFX1 DFF_898_Q_reg ( .D(g25234), .SI(g1554), .SE(test_se), .CLK(CK), .Q(
        g1555), .QN() );
  SDFFX1 DFF_899_Q_reg ( .D(g25242), .SI(g1555), .SE(test_se), .CLK(CK), .Q(
        test_so54), .QN() );
  SDFFX1 DFF_900_Q_reg ( .D(g25235), .SI(test_si55), .SE(test_se), .CLK(CK), 
        .Q(g1557), .QN() );
  SDFFX1 DFF_901_Q_reg ( .D(g25243), .SI(g1557), .SE(test_se), .CLK(CK), .Q(
        g1558), .QN() );
  SDFFX1 DFF_902_Q_reg ( .D(g25249), .SI(g1558), .SE(test_se), .CLK(CK), .Q(
        g1556), .QN() );
  SDFFX1 DFF_903_Q_reg ( .D(g25244), .SI(g1556), .SE(test_se), .CLK(CK), .Q(
        g1560), .QN() );
  SDFFX1 DFF_904_Q_reg ( .D(g25250), .SI(g1560), .SE(test_se), .CLK(CK), .Q(
        g1561), .QN() );
  SDFFX1 DFF_905_Q_reg ( .D(g25255), .SI(g1561), .SE(test_se), .CLK(CK), .Q(
        g1559), .QN() );
  SDFFX1 DFF_906_Q_reg ( .D(g30279), .SI(g1559), .SE(test_se), .CLK(CK), .Q(
        g1567), .QN() );
  SDFFX1 DFF_907_Q_reg ( .D(g30287), .SI(g1567), .SE(test_se), .CLK(CK), .Q(
        g1570), .QN() );
  SDFFX1 DFF_908_Q_reg ( .D(g30294), .SI(g1570), .SE(test_se), .CLK(CK), .Q(
        g1573), .QN() );
  SDFFX1 DFF_909_Q_reg ( .D(g30651), .SI(g1573), .SE(test_se), .CLK(CK), .Q(
        g1612), .QN() );
  SDFFX1 DFF_910_Q_reg ( .D(g30657), .SI(g1612), .SE(test_se), .CLK(CK), .Q(
        g1615), .QN() );
  SDFFX1 DFF_911_Q_reg ( .D(g30663), .SI(g1615), .SE(test_se), .CLK(CK), .Q(
        g1618), .QN() );
  SDFFX1 DFF_912_Q_reg ( .D(g30683), .SI(g1618), .SE(test_se), .CLK(CK), .Q(
        g1576), .QN() );
  SDFFX1 DFF_913_Q_reg ( .D(g30688), .SI(g1576), .SE(test_se), .CLK(CK), .Q(
        g1579), .QN() );
  SDFFX1 DFF_914_Q_reg ( .D(g30692), .SI(g1579), .SE(test_se), .CLK(CK), .Q(
        g1582), .QN() );
  SDFFX1 DFF_915_Q_reg ( .D(g30658), .SI(g1582), .SE(test_se), .CLK(CK), .Q(
        test_so55), .QN() );
  SDFFX1 DFF_916_Q_reg ( .D(g30664), .SI(test_si56), .SE(test_se), .CLK(CK), 
        .Q(g1624), .QN() );
  SDFFX1 DFF_917_Q_reg ( .D(g30671), .SI(g1624), .SE(test_se), .CLK(CK), .Q(
        g1627), .QN() );
  SDFFX1 DFF_918_Q_reg ( .D(g30295), .SI(g1627), .SE(test_se), .CLK(CK), .Q(
        g1585), .QN() );
  SDFFX1 DFF_919_Q_reg ( .D(g30299), .SI(g1585), .SE(test_se), .CLK(CK), .Q(
        g1588), .QN() );
  SDFFX1 DFF_920_Q_reg ( .D(g30302), .SI(g1588), .SE(test_se), .CLK(CK), .Q(
        g1591), .QN() );
  SDFFX1 DFF_921_Q_reg ( .D(g30266), .SI(g1591), .SE(test_se), .CLK(CK), .Q(
        g1630), .QN() );
  SDFFX1 DFF_922_Q_reg ( .D(g30272), .SI(g1630), .SE(test_se), .CLK(CK), .Q(
        g1633), .QN() );
  SDFFX1 DFF_923_Q_reg ( .D(g30280), .SI(g1633), .SE(test_se), .CLK(CK), .Q(
        g1636), .QN() );
  SDFFX1 DFF_924_Q_reg ( .D(g30250), .SI(g1636), .SE(test_se), .CLK(CK), .Q(
        g1594), .QN() );
  SDFFX1 DFF_925_Q_reg ( .D(g30252), .SI(g1594), .SE(test_se), .CLK(CK), .Q(
        g1597), .QN() );
  SDFFX1 DFF_926_Q_reg ( .D(g30255), .SI(g1597), .SE(test_se), .CLK(CK), .Q(
        g1600), .QN() );
  SDFFX1 DFF_927_Q_reg ( .D(g30273), .SI(g1600), .SE(test_se), .CLK(CK), .Q(
        g1639), .QN() );
  SDFFX1 DFF_928_Q_reg ( .D(g30281), .SI(g1639), .SE(test_se), .CLK(CK), .Q(
        g1642), .QN() );
  SDFFX1 DFF_929_Q_reg ( .D(g30288), .SI(g1642), .SE(test_se), .CLK(CK), .Q(
        g1645), .QN() );
  SDFFX1 DFF_930_Q_reg ( .D(g30644), .SI(g1645), .SE(test_se), .CLK(CK), .Q(
        g1603), .QN() );
  SDFFX1 DFF_931_Q_reg ( .D(g30650), .SI(g1603), .SE(test_se), .CLK(CK), .Q(
        test_so56), .QN() );
  SDFFX1 DFF_932_Q_reg ( .D(g30656), .SI(test_si57), .SE(test_se), .CLK(CK), 
        .Q(g1609), .QN() );
  SDFFX1 DFF_933_Q_reg ( .D(g30678), .SI(g1609), .SE(test_se), .CLK(CK), .Q(
        g1648), .QN() );
  SDFFX1 DFF_934_Q_reg ( .D(g30684), .SI(g1648), .SE(test_se), .CLK(CK), .Q(
        g1651), .QN() );
  SDFFX1 DFF_935_Q_reg ( .D(g30689), .SI(g1651), .SE(test_se), .CLK(CK), .Q(
        g1654), .QN() );
  SDFFX1 DFF_936_Q_reg ( .D(g25056), .SI(g1654), .SE(test_se), .CLK(CK), .Q(
        g1466), .QN() );
  SDFFX1 DFF_937_Q_reg ( .D(g25938), .SI(g1466), .SE(test_se), .CLK(CK), .Q(
        g1462), .QN() );
  SDFFX1 DFF_938_Q_reg ( .D(g26531), .SI(g1462), .SE(test_se), .CLK(CK), .Q(
        g1457), .QN() );
  SDFFX1 DFF_939_Q_reg ( .D(g27129), .SI(g1457), .SE(test_se), .CLK(CK), .Q(
        g1453), .QN() );
  SDFFX1 DFF_940_Q_reg ( .D(g27612), .SI(g1453), .SE(test_se), .CLK(CK), .Q(
        g1448), .QN() );
  SDFFX1 DFF_941_Q_reg ( .D(g28147), .SI(g1448), .SE(test_se), .CLK(CK), .Q(
        g1444), .QN() );
  SDFFX1 DFF_942_Q_reg ( .D(g28636), .SI(g1444), .SE(test_se), .CLK(CK), .Q(
        g1439), .QN() );
  SDFFX1 DFF_943_Q_reg ( .D(g29111), .SI(g1439), .SE(test_se), .CLK(CK), .Q(
        g1435), .QN() );
  SDFFX1 DFF_944_Q_reg ( .D(g29355), .SI(g1435), .SE(test_se), .CLK(CK), .Q(
        g1430), .QN() );
  SDFFX1 DFF_945_Q_reg ( .D(g29581), .SI(g1430), .SE(test_se), .CLK(CK), .Q(
        g1426), .QN() );
  SDFFX1 DFF_946_Q_reg ( .D(g13110), .SI(g1426), .SE(test_se), .CLK(CK), .Q(
        g1562), .QN() );
  SDFFX1 DFF_947_Q_reg ( .D(g1562), .SI(g1562), .SE(test_se), .CLK(CK), .Q(
        g5612), .QN() );
  SDFFX1 DFF_948_Q_reg ( .D(g5612), .SI(test_si58), .SE(test_se), .CLK(CK), 
        .Q(g1563), .QN() );
  SDFFX1 DFF_949_Q_reg ( .D(n4650), .SI(g1563), .SE(test_se), .CLK(CK), .Q(
        g1657), .QN(n4518) );
  SDFFX1 DFF_952_Q_reg ( .D(g5612), .SI(g1782), .SE(test_se), .CLK(CK), .Q(
        g1690), .QN(n4386) );
  SDFFX1 DFF_953_Q_reg ( .D(g27264), .SI(g1690), .SE(test_se), .CLK(CK), .Q(
        g1735), .QN() );
  SDFFX1 DFF_954_Q_reg ( .D(g27274), .SI(g1735), .SE(test_se), .CLK(CK), .Q(
        g1724), .QN() );
  SDFFX1 DFF_955_Q_reg ( .D(g27287), .SI(g1724), .SE(test_se), .CLK(CK), .Q(
        g1727), .QN() );
  SDFFX1 DFF_956_Q_reg ( .D(g27275), .SI(g1727), .SE(test_se), .CLK(CK), .Q(
        g1750), .QN() );
  SDFFX1 DFF_957_Q_reg ( .D(g27288), .SI(g1750), .SE(test_se), .CLK(CK), .Q(
        g1739), .QN() );
  SDFFX1 DFF_958_Q_reg ( .D(g27302), .SI(g1739), .SE(test_se), .CLK(CK), .Q(
        g1742), .QN() );
  SDFFX1 DFF_959_Q_reg ( .D(g27289), .SI(g1742), .SE(test_se), .CLK(CK), .Q(
        g1765), .QN() );
  SDFFX1 DFF_960_Q_reg ( .D(g27303), .SI(g1765), .SE(test_se), .CLK(CK), .Q(
        g1754), .QN() );
  SDFFX1 DFF_961_Q_reg ( .D(g27317), .SI(g1754), .SE(test_se), .CLK(CK), .Q(
        g1757), .QN() );
  SDFFX1 DFF_962_Q_reg ( .D(g27304), .SI(g1757), .SE(test_se), .CLK(CK), .Q(
        g1779), .QN() );
  SDFFX1 DFF_963_Q_reg ( .D(g27318), .SI(g1779), .SE(test_se), .CLK(CK), .Q(
        test_so58), .QN() );
  SDFFX1 DFF_964_Q_reg ( .D(g27330), .SI(test_si59), .SE(test_se), .CLK(CK), 
        .Q(g1772), .QN() );
  SDFFX1 DFF_965_Q_reg ( .D(g28749), .SI(g1772), .SE(test_se), .CLK(CK), .Q(
        g1789), .QN() );
  SDFFX1 DFF_966_Q_reg ( .D(g28760), .SI(g1789), .SE(test_se), .CLK(CK), .Q(
        g1792), .QN() );
  SDFFX1 DFF_967_Q_reg ( .D(g28771), .SI(g1792), .SE(test_se), .CLK(CK), .Q(
        g1795), .QN() );
  SDFFX1 DFF_968_Q_reg ( .D(g29205), .SI(g1795), .SE(test_se), .CLK(CK), .Q(
        g1798), .QN() );
  SDFFX1 DFF_969_Q_reg ( .D(g29212), .SI(g1798), .SE(test_se), .CLK(CK), .Q(
        g1801), .QN() );
  SDFFX1 DFF_970_Q_reg ( .D(g29218), .SI(g1801), .SE(test_se), .CLK(CK), .Q(
        g1804), .QN() );
  SDFFX1 DFF_971_Q_reg ( .D(g28761), .SI(g1804), .SE(test_se), .CLK(CK), .Q(
        g1808), .QN() );
  SDFFX1 DFF_972_Q_reg ( .D(g28772), .SI(g1808), .SE(test_se), .CLK(CK), .Q(
        g1809), .QN() );
  SDFFX1 DFF_973_Q_reg ( .D(g28778), .SI(g1809), .SE(test_se), .CLK(CK), .Q(
        g1807), .QN() );
  SDFFX1 DFF_974_Q_reg ( .D(g26811), .SI(g1807), .SE(test_se), .CLK(CK), .Q(
        g1810), .QN() );
  SDFFX1 DFF_975_Q_reg ( .D(g26815), .SI(g1810), .SE(test_se), .CLK(CK), .Q(
        g1813), .QN() );
  SDFFX1 DFF_976_Q_reg ( .D(g26820), .SI(g1813), .SE(test_se), .CLK(CK), .Q(
        g1816), .QN() );
  SDFFX1 DFF_977_Q_reg ( .D(g26816), .SI(g1816), .SE(test_se), .CLK(CK), .Q(
        g1819), .QN() );
  SDFFX1 DFF_978_Q_reg ( .D(g26821), .SI(g1819), .SE(test_se), .CLK(CK), .Q(
        g1822), .QN() );
  SDFFX1 DFF_979_Q_reg ( .D(g26824), .SI(g1822), .SE(test_se), .CLK(CK), .Q(
        test_so59), .QN() );
  SDFFX1 DFF_980_Q_reg ( .D(g27764), .SI(test_si60), .SE(test_se), .CLK(CK), 
        .Q(g1829), .QN() );
  SDFFX1 DFF_981_Q_reg ( .D(g27766), .SI(g1829), .SE(test_se), .CLK(CK), .Q(
        g1830), .QN() );
  SDFFX1 DFF_982_Q_reg ( .D(g27768), .SI(g1830), .SE(test_se), .CLK(CK), .Q(
        g1828), .QN() );
  SDFFX1 DFF_983_Q_reg ( .D(g29613), .SI(g1828), .SE(test_se), .CLK(CK), .Q(
        g1693), .QN() );
  SDFFX1 DFF_984_Q_reg ( .D(g29617), .SI(g1693), .SE(test_se), .CLK(CK), .Q(
        g1694), .QN() );
  SDFFX1 DFF_985_Q_reg ( .D(g29620), .SI(g1694), .SE(test_se), .CLK(CK), .Q(
        g1695), .QN() );
  SDFFX1 DFF_986_Q_reg ( .D(g30704), .SI(g1695), .SE(test_se), .CLK(CK), .Q(
        g1696), .QN() );
  SDFFX1 DFF_987_Q_reg ( .D(g30706), .SI(g1696), .SE(test_se), .CLK(CK), .Q(
        g1697), .QN() );
  SDFFX1 DFF_988_Q_reg ( .D(g30708), .SI(g1697), .SE(test_se), .CLK(CK), .Q(
        g1698), .QN() );
  SDFFX1 DFF_989_Q_reg ( .D(g30487), .SI(g1698), .SE(test_se), .CLK(CK), .Q(
        g1699), .QN() );
  SDFFX1 DFF_990_Q_reg ( .D(g30503), .SI(g1699), .SE(test_se), .CLK(CK), .Q(
        g1700), .QN() );
  SDFFX1 DFF_991_Q_reg ( .D(g30338), .SI(g1700), .SE(test_se), .CLK(CK), .Q(
        g1701), .QN() );
  SDFFX1 DFF_992_Q_reg ( .D(g29178), .SI(g1701), .SE(test_se), .CLK(CK), .Q(
        g1703), .QN() );
  SDFFX1 DFF_993_Q_reg ( .D(g29181), .SI(g1703), .SE(test_se), .CLK(CK), .Q(
        g1704), .QN() );
  SDFFX1 DFF_994_Q_reg ( .D(g29184), .SI(g1704), .SE(test_se), .CLK(CK), .Q(
        g1702), .QN() );
  SDFFX1 DFF_995_Q_reg ( .D(g26667), .SI(g1702), .SE(test_se), .CLK(CK), .Q(
        test_so60), .QN() );
  SDFFX1 DFF_996_Q_reg ( .D(g26670), .SI(test_si61), .SE(test_se), .CLK(CK), 
        .Q(g1785), .QN() );
  SDFFX1 DFF_997_Q_reg ( .D(g26675), .SI(g1785), .SE(test_se), .CLK(CK), .Q(
        g1783), .QN() );
  SDFFX1 DFF_998_Q_reg ( .D(n4288), .SI(g1783), .SE(test_se), .CLK(CK), .Q(
        g1831), .QN() );
  SDFFX1 DFF_999_Q_reg ( .D(g1831), .SI(g1831), .SE(test_se), .CLK(CK), .Q(
        n7988), .QN(DFF_999_n1) );
  SDFFX1 DFF_1000_Q_reg ( .D(n4565), .SI(n7988), .SE(test_se), .CLK(CK), .Q(
        g1833), .QN() );
  SDFFX1 DFF_1001_Q_reg ( .D(g1833), .SI(g1833), .SE(test_se), .CLK(CK), .Q(
        n7987), .QN(DFF_1001_n1) );
  SDFFX1 DFF_1002_Q_reg ( .D(n4557), .SI(n7987), .SE(test_se), .CLK(CK), .Q(
        g1835), .QN() );
  SDFFX1 DFF_1003_Q_reg ( .D(g1835), .SI(g1835), .SE(test_se), .CLK(CK), .Q(
        n7986), .QN(DFF_1003_n1) );
  SDFFX1 DFF_1004_Q_reg ( .D(n4326), .SI(n7986), .SE(test_se), .CLK(CK), .Q(
        g1661), .QN() );
  SDFFX1 DFF_1005_Q_reg ( .D(g1661), .SI(g1661), .SE(test_se), .CLK(CK), .Q(
        n7985), .QN(DFF_1005_n1) );
  SDFFX1 DFF_1006_Q_reg ( .D(n4390), .SI(n7985), .SE(test_se), .CLK(CK), .Q(
        g1663), .QN() );
  SDFFX1 DFF_1007_Q_reg ( .D(g1663), .SI(g1663), .SE(test_se), .CLK(CK), .Q(
        n7984), .QN(DFF_1007_n1) );
  SDFFX1 DFF_1008_Q_reg ( .D(n4320), .SI(n7984), .SE(test_se), .CLK(CK), .Q(
        g1665), .QN() );
  SDFFX1 DFF_1009_Q_reg ( .D(g1665), .SI(g1665), .SE(test_se), .CLK(CK), .Q(
        n7983), .QN(DFF_1009_n1) );
  SDFFX1 DFF_1010_Q_reg ( .D(n4374), .SI(n7983), .SE(test_se), .CLK(CK), .Q(
        g1667), .QN() );
  SDFFX1 DFF_1011_Q_reg ( .D(g1667), .SI(g1667), .SE(test_se), .CLK(CK), .Q(
        test_so61), .QN(DFF_1011_n1) );
  SDFFX1 DFF_1012_Q_reg ( .D(n4378), .SI(test_si62), .SE(test_se), .CLK(CK), 
        .Q(g1669), .QN() );
  SDFFX1 DFF_1013_Q_reg ( .D(g1669), .SI(g1669), .SE(test_se), .CLK(CK), .Q(
        n7980), .QN(DFF_1013_n1) );
  SDFFX1 DFF_1014_Q_reg ( .D(g2877), .SI(n7980), .SE(test_se), .CLK(CK), .Q(
        g1671), .QN() );
  SDFFX1 DFF_1015_Q_reg ( .D(g1671), .SI(g1671), .SE(test_se), .CLK(CK), .Q(
        n7979), .QN(n4484) );
  SDFFX1 DFF_1016_Q_reg ( .D(n4284), .SI(n7979), .SE(test_se), .CLK(CK), .Q(
        g1680), .QN(n4488) );
  SDFFX1 DFF_1017_Q_reg ( .D(g28903), .SI(g1680), .SE(test_se), .CLK(CK), .Q(
        g1686), .QN() );
  SDFFX1 DFF_1028_Q_reg ( .D(n4276), .SI(g1686), .SE(test_se), .CLK(CK), .Q(
        n7978), .QN(n4581) );
  SDFFX1 DFF_1029_Q_reg ( .D(g1735), .SI(n7978), .SE(test_se), .CLK(CK), .Q(
        g1723), .QN() );
  SDFFX1 DFF_1030_Q_reg ( .D(g1723), .SI(g1723), .SE(test_se), .CLK(CK), .Q(
        g1730), .QN() );
  SDFFX1 DFF_1031_Q_reg ( .D(g1724), .SI(g1730), .SE(test_se), .CLK(CK), .Q(
        g1731), .QN() );
  SDFFX1 DFF_1032_Q_reg ( .D(g1731), .SI(g1731), .SE(test_se), .CLK(CK), .Q(
        g1732), .QN() );
  SDFFX1 DFF_1033_Q_reg ( .D(g1727), .SI(g1732), .SE(test_se), .CLK(CK), .Q(
        g1733), .QN() );
  SDFFX1 DFF_1034_Q_reg ( .D(g1733), .SI(g1733), .SE(test_se), .CLK(CK), .Q(
        g1734), .QN() );
  SDFFX1 DFF_1035_Q_reg ( .D(g1750), .SI(g1734), .SE(test_se), .CLK(CK), .Q(
        g1738), .QN() );
  SDFFX1 DFF_1036_Q_reg ( .D(g1738), .SI(g1738), .SE(test_se), .CLK(CK), .Q(
        g1745), .QN() );
  SDFFX1 DFF_1037_Q_reg ( .D(g1739), .SI(g1745), .SE(test_se), .CLK(CK), .Q(
        test_so62), .QN() );
  SDFFX1 DFF_1038_Q_reg ( .D(test_so62), .SI(test_si63), .SE(test_se), .CLK(CK), .Q(g1747), .QN() );
  SDFFX1 DFF_1039_Q_reg ( .D(g1742), .SI(g1747), .SE(test_se), .CLK(CK), .Q(
        g1748), .QN() );
  SDFFX1 DFF_1040_Q_reg ( .D(g1748), .SI(g1748), .SE(test_se), .CLK(CK), .Q(
        g1749), .QN() );
  SDFFX1 DFF_1041_Q_reg ( .D(g1765), .SI(g1749), .SE(test_se), .CLK(CK), .Q(
        g1753), .QN() );
  SDFFX1 DFF_1042_Q_reg ( .D(g1753), .SI(g1753), .SE(test_se), .CLK(CK), .Q(
        g1760), .QN() );
  SDFFX1 DFF_1043_Q_reg ( .D(g1754), .SI(g1760), .SE(test_se), .CLK(CK), .Q(
        g1761), .QN() );
  SDFFX1 DFF_1044_Q_reg ( .D(g1761), .SI(g1761), .SE(test_se), .CLK(CK), .Q(
        g1762), .QN() );
  SDFFX1 DFF_1045_Q_reg ( .D(g1757), .SI(g1762), .SE(test_se), .CLK(CK), .Q(
        g1763), .QN() );
  SDFFX1 DFF_1046_Q_reg ( .D(g1763), .SI(g1763), .SE(test_se), .CLK(CK), .Q(
        g1764), .QN() );
  SDFFX1 DFF_1047_Q_reg ( .D(g1779), .SI(g1764), .SE(test_se), .CLK(CK), .Q(
        g1768), .QN() );
  SDFFX1 DFF_1048_Q_reg ( .D(g1768), .SI(g1768), .SE(test_se), .CLK(CK), .Q(
        g1775), .QN() );
  SDFFX1 DFF_1049_Q_reg ( .D(test_so58), .SI(g1775), .SE(test_se), .CLK(CK), 
        .Q(g1776), .QN() );
  SDFFX1 DFF_1050_Q_reg ( .D(g1776), .SI(g1776), .SE(test_se), .CLK(CK), .Q(
        g1777), .QN() );
  SDFFX1 DFF_1051_Q_reg ( .D(g1772), .SI(g1777), .SE(test_se), .CLK(CK), .Q(
        g1778), .QN() );
  SDFFX1 DFF_1052_Q_reg ( .D(g1778), .SI(g1778), .SE(test_se), .CLK(CK), .Q(
        g1705), .QN() );
  SDFFX1 DFF_1053_Q_reg ( .D(n4598), .SI(g1705), .SE(test_se), .CLK(CK), .Q(
        g5695), .QN() );
  SDFFX1 DFF_1054_Q_reg ( .D(g5695), .SI(test_si64), .SE(test_se), .CLK(CK), 
        .Q(g5738), .QN() );
  SDFFX1 DFF_1055_Q_reg ( .D(g5738), .SI(g5738), .SE(test_se), .CLK(CK), .Q(
        g1718), .QN() );
  SDFFX1 DFF_1056_Q_reg ( .D(n4598), .SI(g1718), .SE(test_se), .CLK(CK), .Q(
        g1925), .QN(n4296) );
  SDFFX1 DFF_1057_Q_reg ( .D(g7052), .SI(g1925), .SE(test_se), .CLK(CK), .Q(
        g1931), .QN(n4315) );
  SDFFX1 DFF_1058_Q_reg ( .D(n4614), .SI(g1931), .SE(test_se), .CLK(CK), .Q(
        g1930), .QN(n4366) );
  SDFFX1 DFF_1059_Q_reg ( .D(g21845), .SI(g1930), .SE(test_se), .CLK(CK), .Q(
        g1934), .QN() );
  SDFFX1 DFF_1060_Q_reg ( .D(g18743), .SI(g1934), .SE(test_se), .CLK(CK), .Q(
        g1937), .QN(n4311) );
  SDFFX1 DFF_1061_Q_reg ( .D(g18794), .SI(g1937), .SE(test_se), .CLK(CK), .Q(
        g1890), .QN(n4297) );
  SDFFX1 DFF_1062_Q_reg ( .D(g12524), .SI(g1890), .SE(test_se), .CLK(CK), .Q(
        g1893), .QN() );
  SDFFX1 DFF_1063_Q_reg ( .D(g1893), .SI(g1893), .SE(test_se), .CLK(CK), .Q(
        g1903), .QN() );
  SDFFX1 DFF_1064_Q_reg ( .D(g1903), .SI(g1903), .SE(test_se), .CLK(CK), .Q(
        g1904), .QN() );
  SDFFX1 DFF_1065_Q_reg ( .D(g1836), .SI(g1904), .SE(test_se), .CLK(CK), .Q(
        g1944), .QN() );
  SDFFX1 DFF_1066_Q_reg ( .D(g1944), .SI(g1944), .SE(test_se), .CLK(CK), .Q(
        g1949), .QN() );
  SDFFX1 DFF_1067_Q_reg ( .D(test_so65), .SI(g1949), .SE(test_se), .CLK(CK), 
        .Q(g1950), .QN() );
  SDFFX1 DFF_1068_Q_reg ( .D(g1950), .SI(g1950), .SE(test_se), .CLK(CK), .Q(
        g1951), .QN() );
  SDFFX1 DFF_1069_Q_reg ( .D(g1842), .SI(g1951), .SE(test_se), .CLK(CK), .Q(
        test_so64), .QN() );
  SDFFX1 DFF_1070_Q_reg ( .D(test_so64), .SI(test_si65), .SE(test_se), .CLK(CK), .Q(g1953), .QN() );
  SDFFX1 DFF_1071_Q_reg ( .D(g1846), .SI(g1953), .SE(test_se), .CLK(CK), .Q(
        g1954), .QN() );
  SDFFX1 DFF_1072_Q_reg ( .D(g1954), .SI(g1954), .SE(test_se), .CLK(CK), .Q(
        g1945), .QN() );
  SDFFX1 DFF_1073_Q_reg ( .D(g1849), .SI(g1945), .SE(test_se), .CLK(CK), .Q(
        g1946), .QN() );
  SDFFX1 DFF_1074_Q_reg ( .D(g1946), .SI(g1946), .SE(test_se), .CLK(CK), .Q(
        g1947), .QN() );
  SDFFX1 DFF_1075_Q_reg ( .D(g1852), .SI(g1947), .SE(test_se), .CLK(CK), .Q(
        g1948), .QN() );
  SDFFX1 DFF_1076_Q_reg ( .D(g1948), .SI(g1948), .SE(test_se), .CLK(CK), .Q(
        g1870), .QN() );
  SDFFX1 DFF_1077_Q_reg ( .D(n4650), .SI(g1870), .SE(test_se), .CLK(CK), .Q(
        g8012), .QN(n4458) );
  SDFFX1 DFF_1078_Q_reg ( .D(g8012), .SI(g8012), .SE(test_se), .CLK(CK), .Q(
        g8082), .QN(n4457) );
  SDFFX1 DFF_1079_Q_reg ( .D(g8082), .SI(g8082), .SE(test_se), .CLK(CK), .Q(
        g1866), .QN(n4464) );
  SDFFX1 DFF_1080_Q_reg ( .D(g23097), .SI(g1866), .SE(test_se), .CLK(CK), .Q(
        g1867), .QN() );
  SDFFX1 DFF_1081_Q_reg ( .D(g23124), .SI(g1867), .SE(test_se), .CLK(CK), .Q(
        g1868), .QN() );
  SDFFX1 DFF_1082_Q_reg ( .D(g23137), .SI(g1868), .SE(test_se), .CLK(CK), .Q(
        g1869), .QN() );
  SDFFX1 DFF_1083_Q_reg ( .D(g23400), .SI(g1869), .SE(test_se), .CLK(CK), .Q(
        g1836), .QN() );
  SDFFX1 DFF_1084_Q_reg ( .D(g23413), .SI(g1836), .SE(test_se), .CLK(CK), .Q(
        test_so65), .QN() );
  SDFFX1 DFF_1085_Q_reg ( .D(g24182), .SI(test_si66), .SE(test_se), .CLK(CK), 
        .Q(g1842), .QN() );
  SDFFX1 DFF_1086_Q_reg ( .D(g24208), .SI(g1842), .SE(test_se), .CLK(CK), .Q(
        g1858), .QN() );
  SDFFX1 DFF_1087_Q_reg ( .D(g24219), .SI(g1858), .SE(test_se), .CLK(CK), .Q(
        g1859), .QN() );
  SDFFX1 DFF_1088_Q_reg ( .D(g24231), .SI(g1859), .SE(test_se), .CLK(CK), .Q(
        g1860), .QN() );
  SDFFX1 DFF_1089_Q_reg ( .D(g23123), .SI(g1860), .SE(test_se), .CLK(CK), .Q(
        g1861), .QN() );
  SDFFX1 DFF_1090_Q_reg ( .D(g23030), .SI(g1861), .SE(test_se), .CLK(CK), .Q(
        g1865), .QN() );
  SDFFX1 DFF_1091_Q_reg ( .D(g23058), .SI(g1865), .SE(test_se), .CLK(CK), .Q(
        g1845), .QN() );
  SDFFX1 DFF_1092_Q_reg ( .D(g24218), .SI(g1845), .SE(test_se), .CLK(CK), .Q(
        g1846), .QN() );
  SDFFX1 DFF_1093_Q_reg ( .D(g24230), .SI(g1846), .SE(test_se), .CLK(CK), .Q(
        g1849), .QN() );
  SDFFX1 DFF_1094_Q_reg ( .D(g24243), .SI(g1849), .SE(test_se), .CLK(CK), .Q(
        g1852), .QN() );
  SDFFX1 DFF_1095_Q_reg ( .D(g12482), .SI(g1852), .SE(test_se), .CLK(CK), .Q(
        g1908), .QN() );
  SDFFX1 DFF_1096_Q_reg ( .D(g1908), .SI(g1908), .SE(test_se), .CLK(CK), .Q(
        g1915), .QN() );
  SDFFX1 DFF_1097_Q_reg ( .D(g1915), .SI(g1915), .SE(test_se), .CLK(CK), .Q(
        g1922), .QN() );
  SDFFX1 DFF_1098_Q_reg ( .D(g13164), .SI(g1922), .SE(test_se), .CLK(CK), .Q(
        g1923), .QN() );
  SDFFX1 DFF_1099_Q_reg ( .D(g1923), .SI(g1923), .SE(test_se), .CLK(CK), .Q(
        test_so66), .QN(DFF_1099_n1) );
  SDFFX1 DFF_1100_Q_reg ( .D(n1818), .SI(test_si67), .SE(test_se), .CLK(CK), 
        .Q(n7971), .QN(DFF_1100_n1) );
  SDFFX1 DFF_1101_Q_reg ( .D(g13135), .SI(n7971), .SE(test_se), .CLK(CK), .Q(
        g1929), .QN() );
  SDFFX1 DFF_1102_Q_reg ( .D(g1929), .SI(g1929), .SE(test_se), .CLK(CK), .Q(
        g1880), .QN(n4545) );
  SDFFX1 DFF_1103_Q_reg ( .D(g13182), .SI(g1880), .SE(test_se), .CLK(CK), .Q(
        g1938), .QN() );
  SDFFX1 DFF_1104_Q_reg ( .D(g1938), .SI(g1938), .SE(test_se), .CLK(CK), .Q(
        g1939), .QN() );
  SDFFX1 DFF_1105_Q_reg ( .D(g27290), .SI(g1939), .SE(test_se), .CLK(CK), .Q(
        g1956), .QN() );
  SDFFX1 DFF_1106_Q_reg ( .D(g27305), .SI(g1956), .SE(test_se), .CLK(CK), .Q(
        g1957), .QN() );
  SDFFX1 DFF_1107_Q_reg ( .D(g27319), .SI(g1957), .SE(test_se), .CLK(CK), .Q(
        g1955), .QN() );
  SDFFX1 DFF_1108_Q_reg ( .D(g27306), .SI(g1955), .SE(test_se), .CLK(CK), .Q(
        g1959), .QN() );
  SDFFX1 DFF_1109_Q_reg ( .D(g27320), .SI(g1959), .SE(test_se), .CLK(CK), .Q(
        g1960), .QN() );
  SDFFX1 DFF_1110_Q_reg ( .D(g27331), .SI(g1960), .SE(test_se), .CLK(CK), .Q(
        g1958), .QN() );
  SDFFX1 DFF_1111_Q_reg ( .D(g27321), .SI(g1958), .SE(test_se), .CLK(CK), .Q(
        g1962), .QN() );
  SDFFX1 DFF_1112_Q_reg ( .D(g27332), .SI(g1962), .SE(test_se), .CLK(CK), .Q(
        g1963), .QN() );
  SDFFX1 DFF_1113_Q_reg ( .D(g27340), .SI(g1963), .SE(test_se), .CLK(CK), .Q(
        g1961), .QN() );
  SDFFX1 DFF_1114_Q_reg ( .D(g27333), .SI(g1961), .SE(test_se), .CLK(CK), .Q(
        test_so67), .QN() );
  SDFFX1 DFF_1115_Q_reg ( .D(g27341), .SI(test_si68), .SE(test_se), .CLK(CK), 
        .Q(g1966), .QN() );
  SDFFX1 DFF_1116_Q_reg ( .D(g27346), .SI(g1966), .SE(test_se), .CLK(CK), .Q(
        g1964), .QN() );
  SDFFX1 DFF_1117_Q_reg ( .D(g24513), .SI(g1964), .SE(test_se), .CLK(CK), .Q(
        g1967), .QN() );
  SDFFX1 DFF_1118_Q_reg ( .D(g24524), .SI(g1967), .SE(test_se), .CLK(CK), .Q(
        g1970), .QN() );
  SDFFX1 DFF_1119_Q_reg ( .D(g24534), .SI(g1970), .SE(test_se), .CLK(CK), .Q(
        g1973), .QN() );
  SDFFX1 DFF_1120_Q_reg ( .D(g24525), .SI(g1973), .SE(test_se), .CLK(CK), .Q(
        g1976), .QN() );
  SDFFX1 DFF_1121_Q_reg ( .D(g24535), .SI(g1976), .SE(test_se), .CLK(CK), .Q(
        g1979), .QN() );
  SDFFX1 DFF_1122_Q_reg ( .D(g24545), .SI(g1979), .SE(test_se), .CLK(CK), .Q(
        g1982), .QN() );
  SDFFX1 DFF_1123_Q_reg ( .D(g28357), .SI(g1982), .SE(test_se), .CLK(CK), .Q(
        g1994), .QN() );
  SDFFX1 DFF_1124_Q_reg ( .D(g28362), .SI(g1994), .SE(test_se), .CLK(CK), .Q(
        g1997), .QN() );
  SDFFX1 DFF_1125_Q_reg ( .D(g28366), .SI(g1997), .SE(test_se), .CLK(CK), .Q(
        g2000), .QN() );
  SDFFX1 DFF_1126_Q_reg ( .D(g28352), .SI(g2000), .SE(test_se), .CLK(CK), .Q(
        g1985), .QN() );
  SDFFX1 DFF_1127_Q_reg ( .D(g28356), .SI(g1985), .SE(test_se), .CLK(CK), .Q(
        g1988), .QN() );
  SDFFX1 DFF_1128_Q_reg ( .D(g28361), .SI(g1988), .SE(test_se), .CLK(CK), .Q(
        g1991), .QN() );
  SDFFX1 DFF_1129_Q_reg ( .D(g26559), .SI(g1991), .SE(test_se), .CLK(CK), .Q(
        test_so68), .QN() );
  SDFFX1 DFF_1130_Q_reg ( .D(g26573), .SI(test_si69), .SE(test_se), .CLK(CK), 
        .Q(g1874), .QN() );
  SDFFX1 DFF_1131_Q_reg ( .D(g26592), .SI(g1874), .SE(test_se), .CLK(CK), .Q(
        g1877), .QN() );
  SDFFX1 DFF_1132_Q_reg ( .D(g1880), .SI(g1877), .SE(test_se), .CLK(CK), .Q(
        g1886), .QN(n4493) );
  SDFFX1 DFF_1133_Q_reg ( .D(g22651), .SI(g1886), .SE(test_se), .CLK(CK), .Q(
        n7968), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(g28990), .SI(n7968), .SE(test_se), .CLK(CK), .Q(
        g16399), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(g16399), .SI(g16399), .SE(test_se), .CLK(CK), .Q(
        g1905), .QN() );
  SDFFX1 DFF_1144_Q_reg ( .D(DFF_999_n1), .SI(g1905), .SE(test_se), .CLK(CK), 
        .Q(n7967), .QN(DFF_1144_n1) );
  SDFFX1 DFF_1145_Q_reg ( .D(DFF_1001_n1), .SI(n7967), .SE(test_se), .CLK(CK), 
        .Q(n7966), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(DFF_1003_n1), .SI(n7966), .SE(test_se), .CLK(CK), 
        .Q(n7965), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(DFF_1005_n1), .SI(n7965), .SE(test_se), .CLK(CK), 
        .Q(n7964), .QN(DFF_1147_n1) );
  SDFFX1 DFF_1148_Q_reg ( .D(DFF_1007_n1), .SI(n7964), .SE(test_se), .CLK(CK), 
        .Q(n7963), .QN(DFF_1148_n1) );
  SDFFX1 DFF_1149_Q_reg ( .D(DFF_1009_n1), .SI(n7963), .SE(test_se), .CLK(CK), 
        .Q(n7962), .QN(DFF_1149_n1) );
  SDFFX1 DFF_1150_Q_reg ( .D(DFF_1011_n1), .SI(n7962), .SE(test_se), .CLK(CK), 
        .Q(g1916), .QN() );
  SDFFX1 DFF_1151_Q_reg ( .D(DFF_1013_n1), .SI(g1916), .SE(test_se), .CLK(CK), 
        .Q(g1917), .QN() );
  SDFFX1 DFF_1152_Q_reg ( .D(g24083), .SI(g1917), .SE(test_se), .CLK(CK), .Q(
        test_so69), .QN(n4491) );
  SDFFX1 DFF_1153_Q_reg ( .D(n4484), .SI(test_si70), .SE(test_se), .CLK(CK), 
        .Q(n7960), .QN(DFF_1153_n1) );
  SDFFX1 DFF_1155_Q_reg ( .D(g7229), .SI(g7229), .SE(test_se), .CLK(CK), .Q(
        g7357), .QN(n4357) );
  SDFFX1 DFF_1156_Q_reg ( .D(g7357), .SI(g7357), .SE(test_se), .CLK(CK), .Q(
        g2009), .QN(n4293) );
  SDFFX1 DFF_1157_Q_reg ( .D(g16692), .SI(g2009), .SE(test_se), .CLK(CK), .Q(
        g2010), .QN() );
  SDFFX1 DFF_1158_Q_reg ( .D(g20353), .SI(g2010), .SE(test_se), .CLK(CK), .Q(
        g2039), .QN(n4427) );
  SDFFX1 DFF_1159_Q_reg ( .D(g20752), .SI(g2039), .SE(test_se), .CLK(CK), .Q(
        g2020), .QN(n4400) );
  SDFFX1 DFF_1160_Q_reg ( .D(g21972), .SI(g2020), .SE(test_se), .CLK(CK), .Q(
        g2013), .QN(n4474) );
  SDFFX1 DFF_1161_Q_reg ( .D(g23339), .SI(g2013), .SE(test_se), .CLK(CK), .Q(
        g2033), .QN(n4420) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24434), .SI(g2033), .SE(test_se), .CLK(CK), .Q(
        g2026), .QN(n4410) );
  SDFFX1 DFF_1163_Q_reg ( .D(g25194), .SI(g2026), .SE(test_se), .CLK(CK), .Q(
        g2040), .QN(n4399) );
  SDFFX1 DFF_1164_Q_reg ( .D(g26671), .SI(g2040), .SE(test_se), .CLK(CK), .Q(
        g2052), .QN(n4409) );
  SDFFX1 DFF_1165_Q_reg ( .D(g26789), .SI(g2052), .SE(test_se), .CLK(CK), .Q(
        g2046), .QN(n4468) );
  SDFFX1 DFF_1166_Q_reg ( .D(g27682), .SI(g2046), .SE(test_se), .CLK(CK), .Q(
        g2059), .QN(n4473) );
  SDFFX1 DFF_1167_Q_reg ( .D(g27722), .SI(g2059), .SE(test_se), .CLK(CK), .Q(
        test_so70), .QN(n4394) );
  SDFFX1 DFF_1168_Q_reg ( .D(g28325), .SI(test_si71), .SE(test_se), .CLK(CK), 
        .Q(g2072), .QN(n4416) );
  SDFFX1 DFF_1169_Q_reg ( .D(g20899), .SI(g2072), .SE(test_se), .CLK(CK), .Q(
        g2079), .QN() );
  SDFFX1 DFF_1170_Q_reg ( .D(g20915), .SI(g2079), .SE(test_se), .CLK(CK), .Q(
        g2080), .QN() );
  SDFFX1 DFF_1171_Q_reg ( .D(g20934), .SI(g2080), .SE(test_se), .CLK(CK), .Q(
        g2078), .QN() );
  SDFFX1 DFF_1172_Q_reg ( .D(g20916), .SI(g2078), .SE(test_se), .CLK(CK), .Q(
        g2082), .QN() );
  SDFFX1 DFF_1173_Q_reg ( .D(g20935), .SI(g2082), .SE(test_se), .CLK(CK), .Q(
        g2083), .QN() );
  SDFFX1 DFF_1174_Q_reg ( .D(g20953), .SI(g2083), .SE(test_se), .CLK(CK), .Q(
        g2081), .QN() );
  SDFFX1 DFF_1175_Q_reg ( .D(g20936), .SI(g2081), .SE(test_se), .CLK(CK), .Q(
        g2085), .QN() );
  SDFFX1 DFF_1176_Q_reg ( .D(g20954), .SI(g2085), .SE(test_se), .CLK(CK), .Q(
        g2086), .QN() );
  SDFFX1 DFF_1177_Q_reg ( .D(g20977), .SI(g2086), .SE(test_se), .CLK(CK), .Q(
        g2084), .QN() );
  SDFFX1 DFF_1178_Q_reg ( .D(g20955), .SI(g2084), .SE(test_se), .CLK(CK), .Q(
        g2088), .QN() );
  SDFFX1 DFF_1179_Q_reg ( .D(g20978), .SI(g2088), .SE(test_se), .CLK(CK), .Q(
        g2089), .QN() );
  SDFFX1 DFF_1180_Q_reg ( .D(g20999), .SI(g2089), .SE(test_se), .CLK(CK), .Q(
        g2087), .QN() );
  SDFFX1 DFF_1181_Q_reg ( .D(g20979), .SI(g2087), .SE(test_se), .CLK(CK), .Q(
        g2091), .QN() );
  SDFFX1 DFF_1182_Q_reg ( .D(g21000), .SI(g2091), .SE(test_se), .CLK(CK), .Q(
        test_so71), .QN() );
  SDFFX1 DFF_1183_Q_reg ( .D(g21019), .SI(test_si72), .SE(test_se), .CLK(CK), 
        .Q(g2090), .QN() );
  SDFFX1 DFF_1184_Q_reg ( .D(g21001), .SI(g2090), .SE(test_se), .CLK(CK), .Q(
        g2094), .QN() );
  SDFFX1 DFF_1185_Q_reg ( .D(g21020), .SI(g2094), .SE(test_se), .CLK(CK), .Q(
        g2095), .QN() );
  SDFFX1 DFF_1186_Q_reg ( .D(g21039), .SI(g2095), .SE(test_se), .CLK(CK), .Q(
        g2093), .QN() );
  SDFFX1 DFF_1187_Q_reg ( .D(g21021), .SI(g2093), .SE(test_se), .CLK(CK), .Q(
        g2097), .QN() );
  SDFFX1 DFF_1188_Q_reg ( .D(g21040), .SI(g2097), .SE(test_se), .CLK(CK), .Q(
        g2098), .QN() );
  SDFFX1 DFF_1189_Q_reg ( .D(g21054), .SI(g2098), .SE(test_se), .CLK(CK), .Q(
        g2096), .QN() );
  SDFFX1 DFF_1190_Q_reg ( .D(g21041), .SI(g2096), .SE(test_se), .CLK(CK), .Q(
        g2100), .QN() );
  SDFFX1 DFF_1191_Q_reg ( .D(g21055), .SI(g2100), .SE(test_se), .CLK(CK), .Q(
        g2101), .QN() );
  SDFFX1 DFF_1192_Q_reg ( .D(g21071), .SI(g2101), .SE(test_se), .CLK(CK), .Q(
        g2099), .QN() );
  SDFFX1 DFF_1193_Q_reg ( .D(g21056), .SI(g2099), .SE(test_se), .CLK(CK), .Q(
        g2103), .QN() );
  SDFFX1 DFF_1194_Q_reg ( .D(g21072), .SI(g2103), .SE(test_se), .CLK(CK), .Q(
        g2104), .QN() );
  SDFFX1 DFF_1195_Q_reg ( .D(g21080), .SI(g2104), .SE(test_se), .CLK(CK), .Q(
        g2102), .QN() );
  SDFFX1 DFF_1196_Q_reg ( .D(g20900), .SI(g2102), .SE(test_se), .CLK(CK), .Q(
        g2106), .QN() );
  SDFFX1 DFF_1197_Q_reg ( .D(g20917), .SI(g2106), .SE(test_se), .CLK(CK), .Q(
        test_so72), .QN() );
  SDFFX1 DFF_1198_Q_reg ( .D(g20937), .SI(test_si73), .SE(test_se), .CLK(CK), 
        .Q(g2105), .QN() );
  SDFFX1 DFF_1199_Q_reg ( .D(g20980), .SI(g2105), .SE(test_se), .CLK(CK), .Q(
        g2109), .QN() );
  SDFFX1 DFF_1200_Q_reg ( .D(g21002), .SI(g2109), .SE(test_se), .CLK(CK), .Q(
        g2110), .QN() );
  SDFFX1 DFF_1201_Q_reg ( .D(g21022), .SI(g2110), .SE(test_se), .CLK(CK), .Q(
        g2108), .QN() );
  SDFFX1 DFF_1202_Q_reg ( .D(g21003), .SI(g2108), .SE(test_se), .CLK(CK), .Q(
        g2112), .QN() );
  SDFFX1 DFF_1203_Q_reg ( .D(g21023), .SI(g2112), .SE(test_se), .CLK(CK), .Q(
        g2113), .QN() );
  SDFFX1 DFF_1204_Q_reg ( .D(g21042), .SI(g2113), .SE(test_se), .CLK(CK), .Q(
        g2111), .QN() );
  SDFFX1 DFF_1205_Q_reg ( .D(g25268), .SI(g2111), .SE(test_se), .CLK(CK), .Q(
        g2115), .QN() );
  SDFFX1 DFF_1206_Q_reg ( .D(g25271), .SI(g2115), .SE(test_se), .CLK(CK), .Q(
        g2116), .QN() );
  SDFFX1 DFF_1207_Q_reg ( .D(g25279), .SI(g2116), .SE(test_se), .CLK(CK), .Q(
        g2114), .QN() );
  SDFFX1 DFF_1208_Q_reg ( .D(g22249), .SI(g2114), .SE(test_se), .CLK(CK), .Q(
        g2118), .QN() );
  SDFFX1 DFF_1209_Q_reg ( .D(g22267), .SI(g2118), .SE(test_se), .CLK(CK), .Q(
        g2119), .QN() );
  SDFFX1 DFF_1210_Q_reg ( .D(g22280), .SI(g2119), .SE(test_se), .CLK(CK), .Q(
        g2117), .QN() );
  SDFFX1 DFF_1211_Q_reg ( .D(n4650), .SI(g2117), .SE(test_se), .CLK(CK), .Q(
        g2214), .QN(n4324) );
  SDFFX1 DFF_1212_Q_reg ( .D(g6837), .SI(g2214), .SE(test_se), .CLK(CK), .Q(
        g7084), .QN(n4514) );
  SDFFX1 DFF_1213_Q_reg ( .D(n4587), .SI(test_si74), .SE(test_se), .CLK(CK), 
        .Q(g2241), .QN(n4367) );
  SDFFX1 DFF_1214_Q_reg ( .D(g22170), .SI(g2241), .SE(test_se), .CLK(CK), .Q(
        g2206), .QN() );
  SDFFX1 DFF_1215_Q_reg ( .D(g22182), .SI(g2206), .SE(test_se), .CLK(CK), .Q(
        g2207), .QN() );
  SDFFX1 DFF_1216_Q_reg ( .D(g22192), .SI(g2207), .SE(test_se), .CLK(CK), .Q(
        g2205), .QN() );
  SDFFX1 DFF_1217_Q_reg ( .D(g22183), .SI(g2205), .SE(test_se), .CLK(CK), .Q(
        g2209), .QN() );
  SDFFX1 DFF_1218_Q_reg ( .D(g22193), .SI(g2209), .SE(test_se), .CLK(CK), .Q(
        g2210), .QN() );
  SDFFX1 DFF_1219_Q_reg ( .D(g22200), .SI(g2210), .SE(test_se), .CLK(CK), .Q(
        g2208), .QN() );
  SDFFX1 DFF_1220_Q_reg ( .D(g22045), .SI(g2208), .SE(test_se), .CLK(CK), .Q(
        g2218), .QN() );
  SDFFX1 DFF_1221_Q_reg ( .D(g22060), .SI(g2218), .SE(test_se), .CLK(CK), .Q(
        g2219), .QN() );
  SDFFX1 DFF_1222_Q_reg ( .D(g22076), .SI(g2219), .SE(test_se), .CLK(CK), .Q(
        g2217), .QN() );
  SDFFX1 DFF_1223_Q_reg ( .D(g22061), .SI(g2217), .SE(test_se), .CLK(CK), .Q(
        g2221), .QN() );
  SDFFX1 DFF_1224_Q_reg ( .D(g22077), .SI(g2221), .SE(test_se), .CLK(CK), .Q(
        g2222), .QN() );
  SDFFX1 DFF_1225_Q_reg ( .D(g22097), .SI(g2222), .SE(test_se), .CLK(CK), .Q(
        g2220), .QN() );
  SDFFX1 DFF_1226_Q_reg ( .D(g22078), .SI(g2220), .SE(test_se), .CLK(CK), .Q(
        g2224), .QN() );
  SDFFX1 DFF_1227_Q_reg ( .D(g22098), .SI(g2224), .SE(test_se), .CLK(CK), .Q(
        test_so74), .QN() );
  SDFFX1 DFF_1228_Q_reg ( .D(g22115), .SI(test_si75), .SE(test_se), .CLK(CK), 
        .Q(g2223), .QN() );
  SDFFX1 DFF_1229_Q_reg ( .D(g22099), .SI(g2223), .SE(test_se), .CLK(CK), .Q(
        g2227), .QN() );
  SDFFX1 DFF_1230_Q_reg ( .D(g22116), .SI(g2227), .SE(test_se), .CLK(CK), .Q(
        g2228), .QN() );
  SDFFX1 DFF_1231_Q_reg ( .D(g22138), .SI(g2228), .SE(test_se), .CLK(CK), .Q(
        g2226), .QN() );
  SDFFX1 DFF_1232_Q_reg ( .D(g22117), .SI(g2226), .SE(test_se), .CLK(CK), .Q(
        g2230), .QN() );
  SDFFX1 DFF_1233_Q_reg ( .D(g22139), .SI(g2230), .SE(test_se), .CLK(CK), .Q(
        g2231), .QN() );
  SDFFX1 DFF_1234_Q_reg ( .D(g22153), .SI(g2231), .SE(test_se), .CLK(CK), .Q(
        g2229), .QN() );
  SDFFX1 DFF_1235_Q_reg ( .D(g22140), .SI(g2229), .SE(test_se), .CLK(CK), .Q(
        g2233), .QN() );
  SDFFX1 DFF_1236_Q_reg ( .D(g22154), .SI(g2233), .SE(test_se), .CLK(CK), .Q(
        g2234), .QN() );
  SDFFX1 DFF_1237_Q_reg ( .D(g22171), .SI(g2234), .SE(test_se), .CLK(CK), .Q(
        g2232), .QN() );
  SDFFX1 DFF_1238_Q_reg ( .D(g22155), .SI(g2232), .SE(test_se), .CLK(CK), .Q(
        g2236), .QN() );
  SDFFX1 DFF_1239_Q_reg ( .D(g22172), .SI(g2236), .SE(test_se), .CLK(CK), .Q(
        g2237), .QN() );
  SDFFX1 DFF_1240_Q_reg ( .D(g22184), .SI(g2237), .SE(test_se), .CLK(CK), .Q(
        g2235), .QN() );
  SDFFX1 DFF_1241_Q_reg ( .D(g22173), .SI(g2235), .SE(test_se), .CLK(CK), .Q(
        g2239), .QN() );
  SDFFX1 DFF_1242_Q_reg ( .D(g22185), .SI(g2239), .SE(test_se), .CLK(CK), .Q(
        test_so75), .QN() );
  SDFFX1 DFF_1243_Q_reg ( .D(g22194), .SI(test_si76), .SE(test_se), .CLK(CK), 
        .Q(g2238), .QN() );
  SDFFX1 DFF_1244_Q_reg ( .D(g25227), .SI(g2238), .SE(test_se), .CLK(CK), .Q(
        g2245), .QN() );
  SDFFX1 DFF_1245_Q_reg ( .D(g25236), .SI(g2245), .SE(test_se), .CLK(CK), .Q(
        g2246), .QN() );
  SDFFX1 DFF_1246_Q_reg ( .D(g25245), .SI(g2246), .SE(test_se), .CLK(CK), .Q(
        g2244), .QN() );
  SDFFX1 DFF_1247_Q_reg ( .D(g25237), .SI(g2244), .SE(test_se), .CLK(CK), .Q(
        g2248), .QN() );
  SDFFX1 DFF_1248_Q_reg ( .D(g25246), .SI(g2248), .SE(test_se), .CLK(CK), .Q(
        g2249), .QN() );
  SDFFX1 DFF_1249_Q_reg ( .D(g25251), .SI(g2249), .SE(test_se), .CLK(CK), .Q(
        g2247), .QN() );
  SDFFX1 DFF_1250_Q_reg ( .D(g25247), .SI(g2247), .SE(test_se), .CLK(CK), .Q(
        g2251), .QN() );
  SDFFX1 DFF_1251_Q_reg ( .D(g25252), .SI(g2251), .SE(test_se), .CLK(CK), .Q(
        g2252), .QN() );
  SDFFX1 DFF_1252_Q_reg ( .D(g25256), .SI(g2252), .SE(test_se), .CLK(CK), .Q(
        g2250), .QN() );
  SDFFX1 DFF_1253_Q_reg ( .D(g25253), .SI(g2250), .SE(test_se), .CLK(CK), .Q(
        g2254), .QN() );
  SDFFX1 DFF_1254_Q_reg ( .D(g25257), .SI(g2254), .SE(test_se), .CLK(CK), .Q(
        g2255), .QN() );
  SDFFX1 DFF_1255_Q_reg ( .D(g25259), .SI(g2255), .SE(test_se), .CLK(CK), .Q(
        g2253), .QN() );
  SDFFX1 DFF_1256_Q_reg ( .D(g30289), .SI(g2253), .SE(test_se), .CLK(CK), .Q(
        g2261), .QN() );
  SDFFX1 DFF_1257_Q_reg ( .D(g30296), .SI(g2261), .SE(test_se), .CLK(CK), .Q(
        test_so76), .QN() );
  SDFFX1 DFF_1258_Q_reg ( .D(g30300), .SI(test_si77), .SE(test_se), .CLK(CK), 
        .Q(g2267), .QN() );
  SDFFX1 DFF_1259_Q_reg ( .D(g30660), .SI(g2267), .SE(test_se), .CLK(CK), .Q(
        g2306), .QN() );
  SDFFX1 DFF_1260_Q_reg ( .D(g30666), .SI(g2306), .SE(test_se), .CLK(CK), .Q(
        g2309), .QN() );
  SDFFX1 DFF_1261_Q_reg ( .D(g30672), .SI(g2309), .SE(test_se), .CLK(CK), .Q(
        g2312), .QN() );
  SDFFX1 DFF_1262_Q_reg ( .D(g30690), .SI(g2312), .SE(test_se), .CLK(CK), .Q(
        g2270), .QN() );
  SDFFX1 DFF_1263_Q_reg ( .D(g30693), .SI(g2270), .SE(test_se), .CLK(CK), .Q(
        g2273), .QN() );
  SDFFX1 DFF_1264_Q_reg ( .D(g30695), .SI(g2273), .SE(test_se), .CLK(CK), .Q(
        g2276), .QN() );
  SDFFX1 DFF_1265_Q_reg ( .D(g30667), .SI(g2276), .SE(test_se), .CLK(CK), .Q(
        g2315), .QN() );
  SDFFX1 DFF_1266_Q_reg ( .D(g30673), .SI(g2315), .SE(test_se), .CLK(CK), .Q(
        g2318), .QN() );
  SDFFX1 DFF_1267_Q_reg ( .D(g30679), .SI(g2318), .SE(test_se), .CLK(CK), .Q(
        g2321), .QN() );
  SDFFX1 DFF_1268_Q_reg ( .D(g30301), .SI(g2321), .SE(test_se), .CLK(CK), .Q(
        g2279), .QN() );
  SDFFX1 DFF_1269_Q_reg ( .D(g30303), .SI(g2279), .SE(test_se), .CLK(CK), .Q(
        g2282), .QN() );
  SDFFX1 DFF_1270_Q_reg ( .D(g30304), .SI(g2282), .SE(test_se), .CLK(CK), .Q(
        g2285), .QN() );
  SDFFX1 DFF_1271_Q_reg ( .D(g30274), .SI(g2285), .SE(test_se), .CLK(CK), .Q(
        g2324), .QN() );
  SDFFX1 DFF_1272_Q_reg ( .D(g30282), .SI(g2324), .SE(test_se), .CLK(CK), .Q(
        test_so77), .QN() );
  SDFFX1 DFF_1273_Q_reg ( .D(g30290), .SI(test_si78), .SE(test_se), .CLK(CK), 
        .Q(g2330), .QN() );
  SDFFX1 DFF_1274_Q_reg ( .D(g30253), .SI(g2330), .SE(test_se), .CLK(CK), .Q(
        g2288), .QN() );
  SDFFX1 DFF_1275_Q_reg ( .D(g30256), .SI(g2288), .SE(test_se), .CLK(CK), .Q(
        g2291), .QN() );
  SDFFX1 DFF_1276_Q_reg ( .D(g30260), .SI(g2291), .SE(test_se), .CLK(CK), .Q(
        g2294), .QN() );
  SDFFX1 DFF_1277_Q_reg ( .D(g30283), .SI(g2294), .SE(test_se), .CLK(CK), .Q(
        g2333), .QN() );
  SDFFX1 DFF_1278_Q_reg ( .D(g30291), .SI(g2333), .SE(test_se), .CLK(CK), .Q(
        g2336), .QN() );
  SDFFX1 DFF_1279_Q_reg ( .D(g30297), .SI(g2336), .SE(test_se), .CLK(CK), .Q(
        g2339), .QN() );
  SDFFX1 DFF_1280_Q_reg ( .D(g30652), .SI(g2339), .SE(test_se), .CLK(CK), .Q(
        g2297), .QN() );
  SDFFX1 DFF_1281_Q_reg ( .D(g30659), .SI(g2297), .SE(test_se), .CLK(CK), .Q(
        g2300), .QN() );
  SDFFX1 DFF_1282_Q_reg ( .D(g30665), .SI(g2300), .SE(test_se), .CLK(CK), .Q(
        g2303), .QN() );
  SDFFX1 DFF_1283_Q_reg ( .D(g30686), .SI(g2303), .SE(test_se), .CLK(CK), .Q(
        g2342), .QN() );
  SDFFX1 DFF_1284_Q_reg ( .D(g30691), .SI(g2342), .SE(test_se), .CLK(CK), .Q(
        g2345), .QN() );
  SDFFX1 DFF_1285_Q_reg ( .D(g30694), .SI(g2345), .SE(test_se), .CLK(CK), .Q(
        g2348), .QN() );
  SDFFX1 DFF_1286_Q_reg ( .D(g25067), .SI(g2348), .SE(test_se), .CLK(CK), .Q(
        g2160), .QN() );
  SDFFX1 DFF_1287_Q_reg ( .D(g25940), .SI(g2160), .SE(test_se), .CLK(CK), .Q(
        test_so78), .QN() );
  SDFFX1 DFF_1288_Q_reg ( .D(g26532), .SI(test_si79), .SE(test_se), .CLK(CK), 
        .Q(g2151), .QN() );
  SDFFX1 DFF_1289_Q_reg ( .D(g27131), .SI(g2151), .SE(test_se), .CLK(CK), .Q(
        g2147), .QN() );
  SDFFX1 DFF_1290_Q_reg ( .D(g27621), .SI(g2147), .SE(test_se), .CLK(CK), .Q(
        g2142), .QN() );
  SDFFX1 DFF_1291_Q_reg ( .D(g28148), .SI(g2142), .SE(test_se), .CLK(CK), .Q(
        g2138), .QN() );
  SDFFX1 DFF_1292_Q_reg ( .D(g28637), .SI(g2138), .SE(test_se), .CLK(CK), .Q(
        g2133), .QN() );
  SDFFX1 DFF_1293_Q_reg ( .D(g29112), .SI(g2133), .SE(test_se), .CLK(CK), .Q(
        g2129), .QN() );
  SDFFX1 DFF_1294_Q_reg ( .D(g29357), .SI(g2129), .SE(test_se), .CLK(CK), .Q(
        g2124), .QN() );
  SDFFX1 DFF_1295_Q_reg ( .D(g29582), .SI(g2124), .SE(test_se), .CLK(CK), .Q(
        g2120), .QN() );
  SDFFX1 DFF_1296_Q_reg ( .D(g13110), .SI(g2120), .SE(test_se), .CLK(CK), .Q(
        g2256), .QN() );
  SDFFX1 DFF_1297_Q_reg ( .D(g2256), .SI(g2256), .SE(test_se), .CLK(CK), .Q(
        g5637), .QN() );
  SDFFX1 DFF_1298_Q_reg ( .D(g5637), .SI(g5637), .SE(test_se), .CLK(CK), .Q(
        g2257), .QN() );
  SDFFX1 DFF_1299_Q_reg ( .D(n4650), .SI(g2257), .SE(test_se), .CLK(CK), .Q(
        g2351), .QN(n4516) );
  SDFFX1 DFF_1302_Q_reg ( .D(g5637), .SI(g2476), .SE(test_se), .CLK(CK), .Q(
        test_so79), .QN(n4385) );
  SDFFX1 DFF_1303_Q_reg ( .D(g27276), .SI(test_si80), .SE(test_se), .CLK(CK), 
        .Q(g2429), .QN() );
  SDFFX1 DFF_1304_Q_reg ( .D(g27291), .SI(g2429), .SE(test_se), .CLK(CK), .Q(
        g2418), .QN() );
  SDFFX1 DFF_1305_Q_reg ( .D(g27307), .SI(g2418), .SE(test_se), .CLK(CK), .Q(
        g2421), .QN() );
  SDFFX1 DFF_1306_Q_reg ( .D(g27292), .SI(g2421), .SE(test_se), .CLK(CK), .Q(
        g2444), .QN() );
  SDFFX1 DFF_1307_Q_reg ( .D(g27308), .SI(g2444), .SE(test_se), .CLK(CK), .Q(
        g2433), .QN() );
  SDFFX1 DFF_1308_Q_reg ( .D(g27322), .SI(g2433), .SE(test_se), .CLK(CK), .Q(
        g2436), .QN() );
  SDFFX1 DFF_1309_Q_reg ( .D(g27309), .SI(g2436), .SE(test_se), .CLK(CK), .Q(
        g2459), .QN() );
  SDFFX1 DFF_1310_Q_reg ( .D(g27323), .SI(g2459), .SE(test_se), .CLK(CK), .Q(
        g2448), .QN() );
  SDFFX1 DFF_1311_Q_reg ( .D(g27334), .SI(g2448), .SE(test_se), .CLK(CK), .Q(
        g2451), .QN() );
  SDFFX1 DFF_1312_Q_reg ( .D(g27324), .SI(g2451), .SE(test_se), .CLK(CK), .Q(
        g2473), .QN() );
  SDFFX1 DFF_1313_Q_reg ( .D(g27335), .SI(g2473), .SE(test_se), .CLK(CK), .Q(
        g2463), .QN() );
  SDFFX1 DFF_1314_Q_reg ( .D(g27342), .SI(g2463), .SE(test_se), .CLK(CK), .Q(
        g2466), .QN() );
  SDFFX1 DFF_1315_Q_reg ( .D(g28763), .SI(g2466), .SE(test_se), .CLK(CK), .Q(
        g2483), .QN() );
  SDFFX1 DFF_1316_Q_reg ( .D(g28773), .SI(g2483), .SE(test_se), .CLK(CK), .Q(
        g2486), .QN() );
  SDFFX1 DFF_1317_Q_reg ( .D(g28782), .SI(g2486), .SE(test_se), .CLK(CK), .Q(
        test_so80), .QN() );
  SDFFX1 DFF_1318_Q_reg ( .D(g29213), .SI(test_si81), .SE(test_se), .CLK(CK), 
        .Q(g2492), .QN() );
  SDFFX1 DFF_1319_Q_reg ( .D(g29221), .SI(g2492), .SE(test_se), .CLK(CK), .Q(
        g2495), .QN() );
  SDFFX1 DFF_1320_Q_reg ( .D(g29226), .SI(g2495), .SE(test_se), .CLK(CK), .Q(
        g2498), .QN() );
  SDFFX1 DFF_1321_Q_reg ( .D(g28774), .SI(g2498), .SE(test_se), .CLK(CK), .Q(
        g2502), .QN() );
  SDFFX1 DFF_1322_Q_reg ( .D(g28783), .SI(g2502), .SE(test_se), .CLK(CK), .Q(
        g2503), .QN() );
  SDFFX1 DFF_1323_Q_reg ( .D(g28788), .SI(g2503), .SE(test_se), .CLK(CK), .Q(
        g2501), .QN() );
  SDFFX1 DFF_1324_Q_reg ( .D(g26817), .SI(g2501), .SE(test_se), .CLK(CK), .Q(
        g2504), .QN() );
  SDFFX1 DFF_1325_Q_reg ( .D(g26822), .SI(g2504), .SE(test_se), .CLK(CK), .Q(
        g2507), .QN() );
  SDFFX1 DFF_1326_Q_reg ( .D(g26825), .SI(g2507), .SE(test_se), .CLK(CK), .Q(
        g2510), .QN() );
  SDFFX1 DFF_1327_Q_reg ( .D(g26823), .SI(g2510), .SE(test_se), .CLK(CK), .Q(
        g2513), .QN() );
  SDFFX1 DFF_1328_Q_reg ( .D(g26826), .SI(g2513), .SE(test_se), .CLK(CK), .Q(
        g2516), .QN() );
  SDFFX1 DFF_1329_Q_reg ( .D(g26827), .SI(g2516), .SE(test_se), .CLK(CK), .Q(
        g2519), .QN() );
  SDFFX1 DFF_1330_Q_reg ( .D(g27767), .SI(g2519), .SE(test_se), .CLK(CK), .Q(
        g2523), .QN() );
  SDFFX1 DFF_1331_Q_reg ( .D(g27769), .SI(g2523), .SE(test_se), .CLK(CK), .Q(
        g2524), .QN() );
  SDFFX1 DFF_1332_Q_reg ( .D(g27771), .SI(g2524), .SE(test_se), .CLK(CK), .Q(
        test_so81), .QN() );
  SDFFX1 DFF_1333_Q_reg ( .D(g29618), .SI(test_si82), .SE(test_se), .CLK(CK), 
        .Q(g2387), .QN() );
  SDFFX1 DFF_1334_Q_reg ( .D(g29621), .SI(g2387), .SE(test_se), .CLK(CK), .Q(
        g2388), .QN() );
  SDFFX1 DFF_1335_Q_reg ( .D(g29623), .SI(g2388), .SE(test_se), .CLK(CK), .Q(
        g2389), .QN() );
  SDFFX1 DFF_1336_Q_reg ( .D(g30707), .SI(g2389), .SE(test_se), .CLK(CK), .Q(
        g2390), .QN() );
  SDFFX1 DFF_1337_Q_reg ( .D(g30709), .SI(g2390), .SE(test_se), .CLK(CK), .Q(
        g2391), .QN() );
  SDFFX1 DFF_1338_Q_reg ( .D(g30566), .SI(g2391), .SE(test_se), .CLK(CK), .Q(
        g2392), .QN() );
  SDFFX1 DFF_1339_Q_reg ( .D(g30505), .SI(g2392), .SE(test_se), .CLK(CK), .Q(
        g2393), .QN() );
  SDFFX1 DFF_1340_Q_reg ( .D(g30341), .SI(g2393), .SE(test_se), .CLK(CK), .Q(
        g2394), .QN() );
  SDFFX1 DFF_1341_Q_reg ( .D(g30356), .SI(g2394), .SE(test_se), .CLK(CK), .Q(
        g2395), .QN() );
  SDFFX1 DFF_1342_Q_reg ( .D(g29182), .SI(g2395), .SE(test_se), .CLK(CK), .Q(
        g2397), .QN() );
  SDFFX1 DFF_1343_Q_reg ( .D(g29185), .SI(g2397), .SE(test_se), .CLK(CK), .Q(
        g2398), .QN() );
  SDFFX1 DFF_1344_Q_reg ( .D(g29187), .SI(g2398), .SE(test_se), .CLK(CK), .Q(
        g2396), .QN() );
  SDFFX1 DFF_1345_Q_reg ( .D(g26672), .SI(g2396), .SE(test_se), .CLK(CK), .Q(
        g2478), .QN() );
  SDFFX1 DFF_1346_Q_reg ( .D(g26676), .SI(g2478), .SE(test_se), .CLK(CK), .Q(
        g2479), .QN() );
  SDFFX1 DFF_1347_Q_reg ( .D(g26025), .SI(g2479), .SE(test_se), .CLK(CK), .Q(
        test_so82), .QN() );
  SDFFX1 DFF_1348_Q_reg ( .D(n4287), .SI(test_si83), .SE(test_se), .CLK(CK), 
        .Q(g2525), .QN() );
  SDFFX1 DFF_1349_Q_reg ( .D(g2525), .SI(g2525), .SE(test_se), .CLK(CK), .Q(
        n7946), .QN(DFF_1349_n1) );
  SDFFX1 DFF_1350_Q_reg ( .D(n4563), .SI(n7946), .SE(test_se), .CLK(CK), .Q(
        g2527), .QN() );
  SDFFX1 DFF_1351_Q_reg ( .D(g2527), .SI(g2527), .SE(test_se), .CLK(CK), .Q(
        n7945), .QN(DFF_1351_n1) );
  SDFFX1 DFF_1352_Q_reg ( .D(n4555), .SI(n7945), .SE(test_se), .CLK(CK), .Q(
        g2529), .QN() );
  SDFFX1 DFF_1353_Q_reg ( .D(g2529), .SI(g2529), .SE(test_se), .CLK(CK), .Q(
        n7944), .QN(DFF_1353_n1) );
  SDFFX1 DFF_1354_Q_reg ( .D(n4325), .SI(n7944), .SE(test_se), .CLK(CK), .Q(
        g2355), .QN() );
  SDFFX1 DFF_1355_Q_reg ( .D(g2355), .SI(g2355), .SE(test_se), .CLK(CK), .Q(
        n7943), .QN(DFF_1355_n1) );
  SDFFX1 DFF_1356_Q_reg ( .D(n4389), .SI(n7943), .SE(test_se), .CLK(CK), .Q(
        g2357), .QN() );
  SDFFX1 DFF_1357_Q_reg ( .D(g2357), .SI(g2357), .SE(test_se), .CLK(CK), .Q(
        n7942), .QN(DFF_1357_n1) );
  SDFFX1 DFF_1358_Q_reg ( .D(n4319), .SI(n7942), .SE(test_se), .CLK(CK), .Q(
        g2359), .QN() );
  SDFFX1 DFF_1359_Q_reg ( .D(g2359), .SI(g2359), .SE(test_se), .CLK(CK), .Q(
        n7941), .QN(DFF_1359_n1) );
  SDFFX1 DFF_1360_Q_reg ( .D(n4373), .SI(n7941), .SE(test_se), .CLK(CK), .Q(
        g2361), .QN() );
  SDFFX1 DFF_1361_Q_reg ( .D(g2361), .SI(g2361), .SE(test_se), .CLK(CK), .Q(
        n7940), .QN(DFF_1361_n1) );
  SDFFX1 DFF_1362_Q_reg ( .D(n4377), .SI(n7940), .SE(test_se), .CLK(CK), .Q(
        test_so83), .QN() );
  SDFFX1 DFF_1363_Q_reg ( .D(test_so83), .SI(test_si84), .SE(test_se), .CLK(CK), .Q(n7938), .QN(DFF_1363_n1) );
  SDFFX1 DFF_1364_Q_reg ( .D(g2878), .SI(n7938), .SE(test_se), .CLK(CK), .Q(
        g2365), .QN() );
  SDFFX1 DFF_1365_Q_reg ( .D(g2365), .SI(g2365), .SE(test_se), .CLK(CK), .Q(
        n7937), .QN(n4483) );
  SDFFX1 DFF_1366_Q_reg ( .D(n4285), .SI(n7937), .SE(test_se), .CLK(CK), .Q(
        g2374), .QN(n4487) );
  SDFFX1 DFF_1367_Q_reg ( .D(g30055), .SI(g2374), .SE(test_se), .CLK(CK), .Q(
        g2380), .QN() );
  SDFFX1 DFF_1378_Q_reg ( .D(n4275), .SI(g2380), .SE(test_se), .CLK(CK), .Q(
        n7936), .QN(DFF_1378_n1) );
  SDFFX1 DFF_1379_Q_reg ( .D(g2429), .SI(n7936), .SE(test_se), .CLK(CK), .Q(
        g2417), .QN() );
  SDFFX1 DFF_1380_Q_reg ( .D(g2417), .SI(g2417), .SE(test_se), .CLK(CK), .Q(
        g2424), .QN() );
  SDFFX1 DFF_1381_Q_reg ( .D(g2418), .SI(g2424), .SE(test_se), .CLK(CK), .Q(
        g2425), .QN() );
  SDFFX1 DFF_1382_Q_reg ( .D(g2425), .SI(g2425), .SE(test_se), .CLK(CK), .Q(
        g2426), .QN() );
  SDFFX1 DFF_1383_Q_reg ( .D(g2421), .SI(g2426), .SE(test_se), .CLK(CK), .Q(
        g2427), .QN() );
  SDFFX1 DFF_1384_Q_reg ( .D(g2427), .SI(g2427), .SE(test_se), .CLK(CK), .Q(
        g2428), .QN() );
  SDFFX1 DFF_1385_Q_reg ( .D(g2444), .SI(g2428), .SE(test_se), .CLK(CK), .Q(
        g2432), .QN() );
  SDFFX1 DFF_1386_Q_reg ( .D(g2432), .SI(g2432), .SE(test_se), .CLK(CK), .Q(
        g2439), .QN() );
  SDFFX1 DFF_1387_Q_reg ( .D(g2433), .SI(g2439), .SE(test_se), .CLK(CK), .Q(
        test_so84), .QN() );
  SDFFX1 DFF_1388_Q_reg ( .D(test_so84), .SI(test_si85), .SE(test_se), .CLK(CK), .Q(g2441), .QN() );
  SDFFX1 DFF_1389_Q_reg ( .D(g2436), .SI(g2441), .SE(test_se), .CLK(CK), .Q(
        g2442), .QN() );
  SDFFX1 DFF_1390_Q_reg ( .D(g2442), .SI(g2442), .SE(test_se), .CLK(CK), .Q(
        g2443), .QN() );
  SDFFX1 DFF_1391_Q_reg ( .D(g2459), .SI(g2443), .SE(test_se), .CLK(CK), .Q(
        g2447), .QN() );
  SDFFX1 DFF_1392_Q_reg ( .D(g2447), .SI(g2447), .SE(test_se), .CLK(CK), .Q(
        g2454), .QN() );
  SDFFX1 DFF_1393_Q_reg ( .D(g2448), .SI(g2454), .SE(test_se), .CLK(CK), .Q(
        g2455), .QN() );
  SDFFX1 DFF_1394_Q_reg ( .D(g2455), .SI(g2455), .SE(test_se), .CLK(CK), .Q(
        g2456), .QN() );
  SDFFX1 DFF_1395_Q_reg ( .D(g2451), .SI(g2456), .SE(test_se), .CLK(CK), .Q(
        g2457), .QN() );
  SDFFX1 DFF_1396_Q_reg ( .D(g2457), .SI(g2457), .SE(test_se), .CLK(CK), .Q(
        g2458), .QN() );
  SDFFX1 DFF_1397_Q_reg ( .D(g2473), .SI(g2458), .SE(test_se), .CLK(CK), .Q(
        g2462), .QN() );
  SDFFX1 DFF_1398_Q_reg ( .D(g2462), .SI(g2462), .SE(test_se), .CLK(CK), .Q(
        g2469), .QN() );
  SDFFX1 DFF_1399_Q_reg ( .D(g2463), .SI(g2469), .SE(test_se), .CLK(CK), .Q(
        g2470), .QN() );
  SDFFX1 DFF_1400_Q_reg ( .D(g2470), .SI(g2470), .SE(test_se), .CLK(CK), .Q(
        g2471), .QN() );
  SDFFX1 DFF_1401_Q_reg ( .D(g2466), .SI(g2471), .SE(test_se), .CLK(CK), .Q(
        g2472), .QN() );
  SDFFX1 DFF_1402_Q_reg ( .D(g2472), .SI(g2472), .SE(test_se), .CLK(CK), .Q(
        test_so85), .QN() );
  SDFFX1 DFF_1403_Q_reg ( .D(n4597), .SI(test_si86), .SE(test_se), .CLK(CK), 
        .Q(g5747), .QN() );
  SDFFX1 DFF_1404_Q_reg ( .D(g5747), .SI(g5747), .SE(test_se), .CLK(CK), .Q(
        g5796), .QN() );
  SDFFX1 DFF_1405_Q_reg ( .D(g5796), .SI(g5796), .SE(test_se), .CLK(CK), .Q(
        g2412), .QN() );
  SDFFX1 DFF_1406_Q_reg ( .D(n4597), .SI(g2412), .SE(test_se), .CLK(CK), .Q(
        g2619), .QN(n4314) );
  SDFFX1 DFF_1407_Q_reg ( .D(g7302), .SI(g2619), .SE(test_se), .CLK(CK), .Q(
        g2625), .QN(n4370) );
  SDFFX1 DFF_1408_Q_reg ( .D(n4602), .SI(g2625), .SE(test_se), .CLK(CK), .Q(
        g2624), .QN(n4299) );
  SDFFX1 DFF_1409_Q_reg ( .D(g21847), .SI(g2624), .SE(test_se), .CLK(CK), .Q(
        g2628), .QN() );
  SDFFX1 DFF_1410_Q_reg ( .D(g18780), .SI(g2628), .SE(test_se), .CLK(CK), .Q(
        g2631), .QN(n4352) );
  SDFFX1 DFF_1411_Q_reg ( .D(g18820), .SI(g2631), .SE(test_se), .CLK(CK), .Q(
        g2584), .QN(n4303) );
  SDFFX1 DFF_1412_Q_reg ( .D(g12539), .SI(g2584), .SE(test_se), .CLK(CK), .Q(
        g2587), .QN() );
  SDFFX1 DFF_1413_Q_reg ( .D(g2587), .SI(g2587), .SE(test_se), .CLK(CK), .Q(
        g2597), .QN() );
  SDFFX1 DFF_1414_Q_reg ( .D(g2597), .SI(g2597), .SE(test_se), .CLK(CK), .Q(
        g2598), .QN() );
  SDFFX1 DFF_1415_Q_reg ( .D(g2530), .SI(g2598), .SE(test_se), .CLK(CK), .Q(
        g2638), .QN() );
  SDFFX1 DFF_1416_Q_reg ( .D(g2638), .SI(g2638), .SE(test_se), .CLK(CK), .Q(
        g2643), .QN() );
  SDFFX1 DFF_1417_Q_reg ( .D(g2533), .SI(g2643), .SE(test_se), .CLK(CK), .Q(
        test_so86), .QN() );
  SDFFX1 DFF_1418_Q_reg ( .D(test_so86), .SI(test_si87), .SE(test_se), .CLK(CK), .Q(g2645), .QN() );
  SDFFX1 DFF_1419_Q_reg ( .D(g2536), .SI(g2645), .SE(test_se), .CLK(CK), .Q(
        g2646), .QN() );
  SDFFX1 DFF_1420_Q_reg ( .D(g2646), .SI(g2646), .SE(test_se), .CLK(CK), .Q(
        g2647), .QN() );
  SDFFX1 DFF_1421_Q_reg ( .D(g2540), .SI(g2647), .SE(test_se), .CLK(CK), .Q(
        g2648), .QN() );
  SDFFX1 DFF_1422_Q_reg ( .D(g2648), .SI(g2648), .SE(test_se), .CLK(CK), .Q(
        g2639), .QN() );
  SDFFX1 DFF_1423_Q_reg ( .D(g2543), .SI(g2639), .SE(test_se), .CLK(CK), .Q(
        g2640), .QN() );
  SDFFX1 DFF_1424_Q_reg ( .D(g2640), .SI(g2640), .SE(test_se), .CLK(CK), .Q(
        g2641), .QN() );
  SDFFX1 DFF_1425_Q_reg ( .D(g2546), .SI(g2641), .SE(test_se), .CLK(CK), .Q(
        g2642), .QN() );
  SDFFX1 DFF_1426_Q_reg ( .D(g2642), .SI(g2642), .SE(test_se), .CLK(CK), .Q(
        g2564), .QN() );
  SDFFX1 DFF_1427_Q_reg ( .D(n4650), .SI(g2564), .SE(test_se), .CLK(CK), .Q(
        g8087), .QN(n4456) );
  SDFFX1 DFF_1428_Q_reg ( .D(g8087), .SI(g8087), .SE(test_se), .CLK(CK), .Q(
        g8167), .QN(n4455) );
  SDFFX1 DFF_1429_Q_reg ( .D(g8167), .SI(g8167), .SE(test_se), .CLK(CK), .Q(
        g2560), .QN(n4463) );
  SDFFX1 DFF_1430_Q_reg ( .D(g23114), .SI(g2560), .SE(test_se), .CLK(CK), .Q(
        g2561), .QN() );
  SDFFX1 DFF_1431_Q_reg ( .D(g23133), .SI(g2561), .SE(test_se), .CLK(CK), .Q(
        g2562), .QN() );
  SDFFX1 DFF_1432_Q_reg ( .D(g21970), .SI(g2562), .SE(test_se), .CLK(CK), .Q(
        test_so87), .QN() );
  SDFFX1 DFF_1433_Q_reg ( .D(g23407), .SI(test_si88), .SE(test_se), .CLK(CK), 
        .Q(g2530), .QN() );
  SDFFX1 DFF_1434_Q_reg ( .D(g23418), .SI(g2530), .SE(test_se), .CLK(CK), .Q(
        g2533), .QN() );
  SDFFX1 DFF_1435_Q_reg ( .D(g24209), .SI(g2533), .SE(test_se), .CLK(CK), .Q(
        g2536), .QN() );
  SDFFX1 DFF_1436_Q_reg ( .D(g24214), .SI(g2536), .SE(test_se), .CLK(CK), .Q(
        g2552), .QN() );
  SDFFX1 DFF_1437_Q_reg ( .D(g24226), .SI(g2552), .SE(test_se), .CLK(CK), .Q(
        g2553), .QN() );
  SDFFX1 DFF_1438_Q_reg ( .D(g24238), .SI(g2553), .SE(test_se), .CLK(CK), .Q(
        g2554), .QN() );
  SDFFX1 DFF_1439_Q_reg ( .D(g23132), .SI(g2554), .SE(test_se), .CLK(CK), .Q(
        g2555), .QN() );
  SDFFX1 DFF_1440_Q_reg ( .D(g23047), .SI(g2555), .SE(test_se), .CLK(CK), .Q(
        g2559), .QN() );
  SDFFX1 DFF_1441_Q_reg ( .D(g23076), .SI(g2559), .SE(test_se), .CLK(CK), .Q(
        g2539), .QN() );
  SDFFX1 DFF_1442_Q_reg ( .D(g24225), .SI(g2539), .SE(test_se), .CLK(CK), .Q(
        g2540), .QN() );
  SDFFX1 DFF_1443_Q_reg ( .D(g24237), .SI(g2540), .SE(test_se), .CLK(CK), .Q(
        g2543), .QN() );
  SDFFX1 DFF_1444_Q_reg ( .D(g24250), .SI(g2543), .SE(test_se), .CLK(CK), .Q(
        g2546), .QN() );
  SDFFX1 DFF_1445_Q_reg ( .D(g12499), .SI(g2546), .SE(test_se), .CLK(CK), .Q(
        g2602), .QN() );
  SDFFX1 DFF_1446_Q_reg ( .D(g2602), .SI(g2602), .SE(test_se), .CLK(CK), .Q(
        g2609), .QN() );
  SDFFX1 DFF_1447_Q_reg ( .D(g2609), .SI(g2609), .SE(test_se), .CLK(CK), .Q(
        test_so88), .QN() );
  SDFFX1 DFF_1448_Q_reg ( .D(g13175), .SI(test_si89), .SE(test_se), .CLK(CK), 
        .Q(g2617), .QN() );
  SDFFX1 DFF_1449_Q_reg ( .D(g2617), .SI(g2617), .SE(test_se), .CLK(CK), .Q(
        n7930), .QN(DFF_1449_n1) );
  SDFFX1 DFF_1450_Q_reg ( .D(g30072), .SI(n7930), .SE(test_se), .CLK(CK), .Q(
        n7929), .QN(DFF_1450_n1) );
  SDFFX1 DFF_1451_Q_reg ( .D(g13143), .SI(n7929), .SE(test_se), .CLK(CK), .Q(
        g2623), .QN() );
  SDFFX1 DFF_1452_Q_reg ( .D(g2623), .SI(g2623), .SE(test_se), .CLK(CK), .Q(
        g2574), .QN(n4543) );
  SDFFX1 DFF_1453_Q_reg ( .D(g13194), .SI(g2574), .SE(test_se), .CLK(CK), .Q(
        g2632), .QN() );
  SDFFX1 DFF_1454_Q_reg ( .D(g2632), .SI(g2632), .SE(test_se), .CLK(CK), .Q(
        g2633), .QN() );
  SDFFX1 DFF_1455_Q_reg ( .D(g27310), .SI(g2633), .SE(test_se), .CLK(CK), .Q(
        g2650), .QN() );
  SDFFX1 DFF_1456_Q_reg ( .D(g27325), .SI(g2650), .SE(test_se), .CLK(CK), .Q(
        g2651), .QN() );
  SDFFX1 DFF_1457_Q_reg ( .D(g27336), .SI(g2651), .SE(test_se), .CLK(CK), .Q(
        g2649), .QN() );
  SDFFX1 DFF_1458_Q_reg ( .D(g27326), .SI(g2649), .SE(test_se), .CLK(CK), .Q(
        g2653), .QN() );
  SDFFX1 DFF_1459_Q_reg ( .D(g27337), .SI(g2653), .SE(test_se), .CLK(CK), .Q(
        g2654), .QN() );
  SDFFX1 DFF_1460_Q_reg ( .D(g27343), .SI(g2654), .SE(test_se), .CLK(CK), .Q(
        g2652), .QN() );
  SDFFX1 DFF_1461_Q_reg ( .D(g27338), .SI(g2652), .SE(test_se), .CLK(CK), .Q(
        g2656), .QN() );
  SDFFX1 DFF_1462_Q_reg ( .D(g27344), .SI(g2656), .SE(test_se), .CLK(CK), .Q(
        test_so89), .QN() );
  SDFFX1 DFF_1463_Q_reg ( .D(g27347), .SI(test_si90), .SE(test_se), .CLK(CK), 
        .Q(g2655), .QN() );
  SDFFX1 DFF_1464_Q_reg ( .D(g27345), .SI(g2655), .SE(test_se), .CLK(CK), .Q(
        g2659), .QN() );
  SDFFX1 DFF_1465_Q_reg ( .D(g27348), .SI(g2659), .SE(test_se), .CLK(CK), .Q(
        g2660), .QN() );
  SDFFX1 DFF_1466_Q_reg ( .D(g27354), .SI(g2660), .SE(test_se), .CLK(CK), .Q(
        g2658), .QN() );
  SDFFX1 DFF_1467_Q_reg ( .D(g24527), .SI(g2658), .SE(test_se), .CLK(CK), .Q(
        g2661), .QN() );
  SDFFX1 DFF_1468_Q_reg ( .D(g24537), .SI(g2661), .SE(test_se), .CLK(CK), .Q(
        g2664), .QN() );
  SDFFX1 DFF_1469_Q_reg ( .D(g24547), .SI(g2664), .SE(test_se), .CLK(CK), .Q(
        g2667), .QN() );
  SDFFX1 DFF_1470_Q_reg ( .D(g24538), .SI(g2667), .SE(test_se), .CLK(CK), .Q(
        g2670), .QN() );
  SDFFX1 DFF_1471_Q_reg ( .D(g24548), .SI(g2670), .SE(test_se), .CLK(CK), .Q(
        g2673), .QN() );
  SDFFX1 DFF_1472_Q_reg ( .D(g24557), .SI(g2673), .SE(test_se), .CLK(CK), .Q(
        g2676), .QN() );
  SDFFX1 DFF_1473_Q_reg ( .D(g28364), .SI(g2676), .SE(test_se), .CLK(CK), .Q(
        g2688), .QN() );
  SDFFX1 DFF_1474_Q_reg ( .D(g28368), .SI(g2688), .SE(test_se), .CLK(CK), .Q(
        g2691), .QN() );
  SDFFX1 DFF_1475_Q_reg ( .D(g28371), .SI(g2691), .SE(test_se), .CLK(CK), .Q(
        g2694), .QN() );
  SDFFX1 DFF_1476_Q_reg ( .D(g28358), .SI(g2694), .SE(test_se), .CLK(CK), .Q(
        g2679), .QN() );
  SDFFX1 DFF_1477_Q_reg ( .D(g28363), .SI(g2679), .SE(test_se), .CLK(CK), .Q(
        test_so90), .QN() );
  SDFFX1 DFF_1478_Q_reg ( .D(g28367), .SI(test_si91), .SE(test_se), .CLK(CK), 
        .Q(g2685), .QN() );
  SDFFX1 DFF_1479_Q_reg ( .D(g26575), .SI(g2685), .SE(test_se), .CLK(CK), .Q(
        g2565), .QN() );
  SDFFX1 DFF_1480_Q_reg ( .D(g26596), .SI(g2565), .SE(test_se), .CLK(CK), .Q(
        g2568), .QN() );
  SDFFX1 DFF_1481_Q_reg ( .D(g26616), .SI(g2568), .SE(test_se), .CLK(CK), .Q(
        g2571), .QN() );
  SDFFX1 DFF_1482_Q_reg ( .D(g2574), .SI(g2571), .SE(test_se), .CLK(CK), .Q(
        g2580), .QN() );
  SDFFX1 DFF_1483_Q_reg ( .D(g22687), .SI(g2580), .SE(test_se), .CLK(CK), .Q(
        n7926), .QN(n4579) );
  SDFFX1 DFF_1492_Q_reg ( .D(g30061), .SI(n7926), .SE(test_se), .CLK(CK), .Q(
        g16437), .QN() );
  SDFFX1 DFF_1493_Q_reg ( .D(g16437), .SI(g16437), .SE(test_se), .CLK(CK), .Q(
        g2599), .QN() );
  SDFFX1 DFF_1494_Q_reg ( .D(DFF_1349_n1), .SI(g2599), .SE(test_se), .CLK(CK), 
        .Q(n7925), .QN(DFF_1494_n1) );
  SDFFX1 DFF_1495_Q_reg ( .D(DFF_1351_n1), .SI(n7925), .SE(test_se), .CLK(CK), 
        .Q(n7924), .QN(DFF_1495_n1) );
  SDFFX1 DFF_1496_Q_reg ( .D(DFF_1353_n1), .SI(n7924), .SE(test_se), .CLK(CK), 
        .Q(n7923), .QN(DFF_1496_n1) );
  SDFFX1 DFF_1497_Q_reg ( .D(DFF_1355_n1), .SI(n7923), .SE(test_se), .CLK(CK), 
        .Q(n7922), .QN(DFF_1497_n1) );
  SDFFX1 DFF_1498_Q_reg ( .D(DFF_1357_n1), .SI(n7922), .SE(test_se), .CLK(CK), 
        .Q(n7921), .QN(DFF_1498_n1) );
  SDFFX1 DFF_1499_Q_reg ( .D(DFF_1359_n1), .SI(n7921), .SE(test_se), .CLK(CK), 
        .Q(n7920), .QN(DFF_1499_n1) );
  SDFFX1 DFF_1500_Q_reg ( .D(DFF_1361_n1), .SI(n7920), .SE(test_se), .CLK(CK), 
        .Q(test_so91), .QN() );
  SDFFX1 DFF_1501_Q_reg ( .D(DFF_1363_n1), .SI(test_si92), .SE(test_se), .CLK(
        CK), .Q(g2611), .QN() );
  SDFFX1 DFF_1502_Q_reg ( .D(g24092), .SI(g2611), .SE(test_se), .CLK(CK), .Q(
        g2612), .QN(n4490) );
  SDFFX1 DFF_1503_Q_reg ( .D(n4483), .SI(g2612), .SE(test_se), .CLK(CK), .Q(
        n7918), .QN(DFF_1503_n1) );
  SDFFX1 DFF_1505_Q_reg ( .D(g7425), .SI(g7425), .SE(test_se), .CLK(CK), .Q(
        g7487), .QN(n4356) );
  SDFFX1 DFF_1506_Q_reg ( .D(g7487), .SI(g7487), .SE(test_se), .CLK(CK), .Q(
        g2703), .QN(n4292) );
  SDFFX1 DFF_1507_Q_reg ( .D(g16718), .SI(g2703), .SE(test_se), .CLK(CK), .Q(
        g2704), .QN() );
  SDFFX1 DFF_1508_Q_reg ( .D(g20375), .SI(g2704), .SE(test_se), .CLK(CK), .Q(
        g2733), .QN(n4426) );
  SDFFX1 DFF_1509_Q_reg ( .D(g20789), .SI(g2733), .SE(test_se), .CLK(CK), .Q(
        g2714), .QN(n4398) );
  SDFFX1 DFF_1510_Q_reg ( .D(g21974), .SI(g2714), .SE(test_se), .CLK(CK), .Q(
        g2707), .QN(n4472) );
  SDFFX1 DFF_1511_Q_reg ( .D(g23348), .SI(g2707), .SE(test_se), .CLK(CK), .Q(
        g2727), .QN(n4419) );
  SDFFX1 DFF_1512_Q_reg ( .D(g24438), .SI(g2727), .SE(test_se), .CLK(CK), .Q(
        g2720), .QN(n4408) );
  SDFFX1 DFF_1513_Q_reg ( .D(g25197), .SI(g2720), .SE(test_se), .CLK(CK), .Q(
        g2734), .QN(n4397) );
  SDFFX1 DFF_1514_Q_reg ( .D(g26677), .SI(g2734), .SE(test_se), .CLK(CK), .Q(
        g2746), .QN(n4407) );
  SDFFX1 DFF_1515_Q_reg ( .D(g26795), .SI(g2746), .SE(test_se), .CLK(CK), .Q(
        test_so92), .QN(n4467) );
  SDFFX1 DFF_1516_Q_reg ( .D(g27243), .SI(test_si93), .SE(test_se), .CLK(CK), 
        .Q(g2753), .QN(n4471) );
  SDFFX1 DFF_1517_Q_reg ( .D(g27724), .SI(g2753), .SE(test_se), .CLK(CK), .Q(
        g2760), .QN(n4393) );
  SDFFX1 DFF_1518_Q_reg ( .D(g28328), .SI(g2760), .SE(test_se), .CLK(CK), .Q(
        g2766), .QN(n4415) );
  SDFFX1 DFF_1519_Q_reg ( .D(g20918), .SI(g2766), .SE(test_se), .CLK(CK), .Q(
        g2773), .QN() );
  SDFFX1 DFF_1520_Q_reg ( .D(g20939), .SI(g2773), .SE(test_se), .CLK(CK), .Q(
        g2774), .QN() );
  SDFFX1 DFF_1521_Q_reg ( .D(g20962), .SI(g2774), .SE(test_se), .CLK(CK), .Q(
        g2772), .QN() );
  SDFFX1 DFF_1522_Q_reg ( .D(g20940), .SI(g2772), .SE(test_se), .CLK(CK), .Q(
        g2776), .QN() );
  SDFFX1 DFF_1523_Q_reg ( .D(g20963), .SI(g2776), .SE(test_se), .CLK(CK), .Q(
        g2777), .QN() );
  SDFFX1 DFF_1524_Q_reg ( .D(g20981), .SI(g2777), .SE(test_se), .CLK(CK), .Q(
        g2775), .QN() );
  SDFFX1 DFF_1525_Q_reg ( .D(g20964), .SI(g2775), .SE(test_se), .CLK(CK), .Q(
        g2779), .QN() );
  SDFFX1 DFF_1526_Q_reg ( .D(g20982), .SI(g2779), .SE(test_se), .CLK(CK), .Q(
        g2780), .QN() );
  SDFFX1 DFF_1527_Q_reg ( .D(g21004), .SI(g2780), .SE(test_se), .CLK(CK), .Q(
        g2778), .QN() );
  SDFFX1 DFF_1528_Q_reg ( .D(g20983), .SI(g2778), .SE(test_se), .CLK(CK), .Q(
        g2782), .QN() );
  SDFFX1 DFF_1529_Q_reg ( .D(g21005), .SI(g2782), .SE(test_se), .CLK(CK), .Q(
        g2783), .QN() );
  SDFFX1 DFF_1530_Q_reg ( .D(g21025), .SI(g2783), .SE(test_se), .CLK(CK), .Q(
        test_so93), .QN() );
  SDFFX1 DFF_1531_Q_reg ( .D(g21006), .SI(test_si94), .SE(test_se), .CLK(CK), 
        .Q(g2785), .QN() );
  SDFFX1 DFF_1532_Q_reg ( .D(g21026), .SI(g2785), .SE(test_se), .CLK(CK), .Q(
        g2786), .QN() );
  SDFFX1 DFF_1533_Q_reg ( .D(g21043), .SI(g2786), .SE(test_se), .CLK(CK), .Q(
        g2784), .QN() );
  SDFFX1 DFF_1534_Q_reg ( .D(g21027), .SI(g2784), .SE(test_se), .CLK(CK), .Q(
        g2788), .QN() );
  SDFFX1 DFF_1535_Q_reg ( .D(g21044), .SI(g2788), .SE(test_se), .CLK(CK), .Q(
        g2789), .QN() );
  SDFFX1 DFF_1536_Q_reg ( .D(g21060), .SI(g2789), .SE(test_se), .CLK(CK), .Q(
        g2787), .QN() );
  SDFFX1 DFF_1537_Q_reg ( .D(g21045), .SI(g2787), .SE(test_se), .CLK(CK), .Q(
        g2791), .QN() );
  SDFFX1 DFF_1538_Q_reg ( .D(g21061), .SI(g2791), .SE(test_se), .CLK(CK), .Q(
        g2792), .QN() );
  SDFFX1 DFF_1539_Q_reg ( .D(g21073), .SI(g2792), .SE(test_se), .CLK(CK), .Q(
        g2790), .QN() );
  SDFFX1 DFF_1540_Q_reg ( .D(g21062), .SI(g2790), .SE(test_se), .CLK(CK), .Q(
        g2794), .QN() );
  SDFFX1 DFF_1541_Q_reg ( .D(g21074), .SI(g2794), .SE(test_se), .CLK(CK), .Q(
        g2795), .QN() );
  SDFFX1 DFF_1542_Q_reg ( .D(g21081), .SI(g2795), .SE(test_se), .CLK(CK), .Q(
        g2793), .QN() );
  SDFFX1 DFF_1543_Q_reg ( .D(g21075), .SI(g2793), .SE(test_se), .CLK(CK), .Q(
        g2797), .QN() );
  SDFFX1 DFF_1544_Q_reg ( .D(g21082), .SI(g2797), .SE(test_se), .CLK(CK), .Q(
        g2798), .QN() );
  SDFFX1 DFF_1545_Q_reg ( .D(g21094), .SI(g2798), .SE(test_se), .CLK(CK), .Q(
        test_so94), .QN() );
  SDFFX1 DFF_1546_Q_reg ( .D(g20919), .SI(test_si95), .SE(test_se), .CLK(CK), 
        .Q(g2800), .QN() );
  SDFFX1 DFF_1547_Q_reg ( .D(g20941), .SI(g2800), .SE(test_se), .CLK(CK), .Q(
        g2801), .QN() );
  SDFFX1 DFF_1548_Q_reg ( .D(g20965), .SI(g2801), .SE(test_se), .CLK(CK), .Q(
        g2799), .QN() );
  SDFFX1 DFF_1549_Q_reg ( .D(g21007), .SI(g2799), .SE(test_se), .CLK(CK), .Q(
        g2803), .QN() );
  SDFFX1 DFF_1550_Q_reg ( .D(g21028), .SI(g2803), .SE(test_se), .CLK(CK), .Q(
        g2804), .QN() );
  SDFFX1 DFF_1551_Q_reg ( .D(g21046), .SI(g2804), .SE(test_se), .CLK(CK), .Q(
        g2802), .QN() );
  SDFFX1 DFF_1552_Q_reg ( .D(g21029), .SI(g2802), .SE(test_se), .CLK(CK), .Q(
        g2806), .QN() );
  SDFFX1 DFF_1553_Q_reg ( .D(g21047), .SI(g2806), .SE(test_se), .CLK(CK), .Q(
        g2807), .QN() );
  SDFFX1 DFF_1554_Q_reg ( .D(g21063), .SI(g2807), .SE(test_se), .CLK(CK), .Q(
        g2805), .QN() );
  SDFFX1 DFF_1555_Q_reg ( .D(g25272), .SI(g2805), .SE(test_se), .CLK(CK), .Q(
        g2809), .QN() );
  SDFFX1 DFF_1556_Q_reg ( .D(g25280), .SI(g2809), .SE(test_se), .CLK(CK), .Q(
        g2810), .QN() );
  SDFFX1 DFF_1557_Q_reg ( .D(g25288), .SI(g2810), .SE(test_se), .CLK(CK), .Q(
        g2808), .QN() );
  SDFFX1 DFF_1558_Q_reg ( .D(g22269), .SI(g2808), .SE(test_se), .CLK(CK), .Q(
        g2812), .QN() );
  SDFFX1 DFF_1559_Q_reg ( .D(g22284), .SI(g2812), .SE(test_se), .CLK(CK), .Q(
        g2813), .QN() );
  SDFFX1 DFF_1560_Q_reg ( .D(g22299), .SI(g2813), .SE(test_se), .CLK(CK), .Q(
        test_so95), .QN() );
  SDFFX1 DFF_1561_Q_reg ( .D(g20877), .SI(test_si96), .SE(test_se), .CLK(CK), 
        .Q(n7913), .QN(DFF_1561_n1) );
  SDFFX1 DFF_1562_Q_reg ( .D(g20884), .SI(n7913), .SE(test_se), .CLK(CK), .Q(
        n7912), .QN(DFF_1562_n1) );
  SDFFX1 DFF_1563_Q_reg ( .D(n4263_Tj_Payload), .SI(n7912), .SE(test_se), .CLK(CK), .Q(
        g3080), .QN() );
  SDFFX1 DFF_1564_Q_reg ( .D(n4269), .SI(g3080), .SE(test_se), .CLK(CK), .Q(
        g3043), .QN() );
  SDFFX1 DFF_1565_Q_reg ( .D(n4268), .SI(g3043), .SE(test_se), .CLK(CK), .Q(
        g3044), .QN() );
  SDFFX1 DFF_1566_Q_reg ( .D(n4267), .SI(g3044), .SE(test_se), .CLK(CK), .Q(
        g3045), .QN() );
  SDFFX1 DFF_1567_Q_reg ( .D(n4266), .SI(g3045), .SE(test_se), .CLK(CK), .Q(
        g3046), .QN() );
  SDFFX1 DFF_1568_Q_reg ( .D(n4265), .SI(g3046), .SE(test_se), .CLK(CK), .Q(
        g3047), .QN() );
  SDFFX1 DFF_1569_Q_reg ( .D(n4272), .SI(g3047), .SE(test_se), .CLK(CK), .Q(
        g3048), .QN() );
  SDFFX1 DFF_1570_Q_reg ( .D(n4271), .SI(g3048), .SE(test_se), .CLK(CK), .Q(
        g3049), .QN() );
  SDFFX1 DFF_1571_Q_reg ( .D(n4270), .SI(g3049), .SE(test_se), .CLK(CK), .Q(
        g3050), .QN() );
  SDFFX1 DFF_1572_Q_reg ( .D(n4259), .SI(g3050), .SE(test_se), .CLK(CK), .Q(
        g3051), .QN() );
  SDFFX1 DFF_1573_Q_reg ( .D(n4236), .SI(g3051), .SE(test_se), .CLK(CK), .Q(
        g3052), .QN() );
  SDFFX1 DFF_1574_Q_reg ( .D(n4239), .SI(g3052), .SE(test_se), .CLK(CK), .Q(
        g3053), .QN() );
  SDFFX1 DFF_1575_Q_reg ( .D(n4237), .SI(g3053), .SE(test_se), .CLK(CK), .Q(
        test_so96), .QN() );
  SDFFX1 DFF_1576_Q_reg ( .D(n4234), .SI(test_si97), .SE(test_se), .CLK(CK), 
        .Q(g3056), .QN() );
  SDFFX1 DFF_1577_Q_reg ( .D(n4233), .SI(g3056), .SE(test_se), .CLK(CK), .Q(
        g3057), .QN() );
  SDFFX1 DFF_1578_Q_reg ( .D(n4238), .SI(g3057), .SE(test_se), .CLK(CK), .Q(
        g3058), .QN() );
  SDFFX1 DFF_1579_Q_reg ( .D(n4235), .SI(g3058), .SE(test_se), .CLK(CK), .Q(
        g3059), .QN() );
  SDFFX1 DFF_1580_Q_reg ( .D(n4240), .SI(g3059), .SE(test_se), .CLK(CK), .Q(
        g3060), .QN() );
  SDFFX1 DFF_1581_Q_reg ( .D(n4232), .SI(g3060), .SE(test_se), .CLK(CK), .Q(
        g3061), .QN() );
  SDFFX1 DFF_1582_Q_reg ( .D(n4245), .SI(g3061), .SE(test_se), .CLK(CK), .Q(
        g3062), .QN() );
  SDFFX1 DFF_1583_Q_reg ( .D(n4248), .SI(g3062), .SE(test_se), .CLK(CK), .Q(
        g3063), .QN() );
  SDFFX1 DFF_1584_Q_reg ( .D(n4246), .SI(g3063), .SE(test_se), .CLK(CK), .Q(
        g3064), .QN() );
  SDFFX1 DFF_1585_Q_reg ( .D(n4243), .SI(g3064), .SE(test_se), .CLK(CK), .Q(
        g3065), .QN() );
  SDFFX1 DFF_1586_Q_reg ( .D(n4242), .SI(g3065), .SE(test_se), .CLK(CK), .Q(
        g3066), .QN() );
  SDFFX1 DFF_1587_Q_reg ( .D(n4247), .SI(g3066), .SE(test_se), .CLK(CK), .Q(
        g3067), .QN() );
  SDFFX1 DFF_1588_Q_reg ( .D(n4244), .SI(g3067), .SE(test_se), .CLK(CK), .Q(
        g3068), .QN() );
  SDFFX1 DFF_1589_Q_reg ( .D(n4249), .SI(g3068), .SE(test_se), .CLK(CK), .Q(
        g3069), .QN() );
  SDFFX1 DFF_1590_Q_reg ( .D(n4241), .SI(g3069), .SE(test_se), .CLK(CK), .Q(
        test_so97), .QN() );
  SDFFX1 DFF_1591_Q_reg ( .D(n4254), .SI(test_si98), .SE(test_se), .CLK(CK), 
        .Q(g3071), .QN() );
  SDFFX1 DFF_1592_Q_reg ( .D(n4257), .SI(g3071), .SE(test_se), .CLK(CK), .Q(
        g3072), .QN() );
  SDFFX1 DFF_1593_Q_reg ( .D(n4255), .SI(g3072), .SE(test_se), .CLK(CK), .Q(
        g3073), .QN() );
  SDFFX1 DFF_1594_Q_reg ( .D(n4252), .SI(g3073), .SE(test_se), .CLK(CK), .Q(
        g3074), .QN() );
  SDFFX1 DFF_1595_Q_reg ( .D(n4251), .SI(g3074), .SE(test_se), .CLK(CK), .Q(
        g3075), .QN() );
  SDFFX1 DFF_1596_Q_reg ( .D(n4256), .SI(g3075), .SE(test_se), .CLK(CK), .Q(
        g3076), .QN() );
  SDFFX1 DFF_1597_Q_reg ( .D(n4253), .SI(g3076), .SE(test_se), .CLK(CK), .Q(
        g3077), .QN() );
  SDFFX1 DFF_1598_Q_reg ( .D(n4258), .SI(g3077), .SE(test_se), .CLK(CK), .Q(
        g3078), .QN() );
  SDFFX1 DFF_1599_Q_reg ( .D(n4250), .SI(g3078), .SE(test_se), .CLK(CK), .Q(
        g2997), .QN() );
  SDFFX1 DFF_1600_Q_reg ( .D(g25265), .SI(g2997), .SE(test_se), .CLK(CK), .Q(
        g2993), .QN() );
  SDFFX1 DFF_1601_Q_reg ( .D(g26048), .SI(g2993), .SE(test_se), .CLK(CK), .Q(
        n7909), .QN(n4354) );
  SDFFX1 DFF_1602_Q_reg ( .D(g23330), .SI(n7909), .SE(test_se), .CLK(CK), .Q(
        g3006), .QN() );
  SDFFX1 DFF_1603_Q_reg ( .D(g24445), .SI(g3006), .SE(test_se), .CLK(CK), .Q(
        g3002), .QN() );
  SDFFX1 DFF_1604_Q_reg ( .D(g25191), .SI(g3002), .SE(test_se), .CLK(CK), .Q(
        g3013), .QN() );
  SDFFX1 DFF_1605_Q_reg ( .D(g26031), .SI(g3013), .SE(test_se), .CLK(CK), .Q(
        test_so98), .QN() );
  SDFFX1 DFF_1606_Q_reg ( .D(g26786), .SI(test_si99), .SE(test_se), .CLK(CK), 
        .Q(g3024), .QN() );
  SDFFX1 DFF_1607_Q_reg ( .D(n4262), .SI(g3024), .SE(test_se), .CLK(CK), .Q(
        g3018), .QN(n4481) );
  SDFFX1 DFF_1608_Q_reg ( .D(g23359), .SI(g3018), .SE(test_se), .CLK(CK), .Q(
        g3028), .QN(n4350) );
  SDFFX1 DFF_1609_Q_reg ( .D(g24446), .SI(g3028), .SE(test_se), .CLK(CK), .Q(
        g3036), .QN(n4480) );
  SDFFX1 DFF_1610_Q_reg ( .D(g25202), .SI(g3036), .SE(test_se), .CLK(CK), .Q(
        g3032), .QN() );
  SDFFX1 DFF_1611_Q_reg ( .D(g3234), .SI(g3032), .SE(test_se), .CLK(CK), .Q(
        g5388), .QN() );
  SDFFX1 DFF_1612_Q_reg ( .D(g5388), .SI(g5388), .SE(test_se), .CLK(CK), .Q(
        n7907), .QN(DFF_1612_n1) );
  SDFFX1 DFF_1613_Q_reg ( .D(g16496), .SI(n7907), .SE(test_se), .CLK(CK), .Q(
        g2987), .QN(n4365) );
  SDFFX1 DFF_1614_Q_reg ( .D(g16824), .SI(g2987), .SE(test_se), .CLK(CK), .Q(
        g8275), .QN() );
  SDFFX1 DFF_1615_Q_reg ( .D(g16844), .SI(g8275), .SE(test_se), .CLK(CK), .Q(
        g8274), .QN() );
  SDFFX1 DFF_1616_Q_reg ( .D(g16853), .SI(g8274), .SE(test_se), .CLK(CK), .Q(
        g8273), .QN(DFF_1616_n1) );
  SDFFX1 DFF_1617_Q_reg ( .D(g16860), .SI(g8273), .SE(test_se), .CLK(CK), .Q(
        g8272), .QN(DFF_1617_n1) );
  SDFFX1 DFF_1618_Q_reg ( .D(g16803), .SI(g8272), .SE(test_se), .CLK(CK), .Q(
        g8268), .QN(DFF_1618_n1) );
  SDFFX1 DFF_1619_Q_reg ( .D(g16835), .SI(g8268), .SE(test_se), .CLK(CK), .Q(
        g8269), .QN() );
  SDFFX1 DFF_1620_Q_reg ( .D(g16851), .SI(g8269), .SE(test_se), .CLK(CK), .Q(
        g8270), .QN() );
  SDFFX1 DFF_1621_Q_reg ( .D(g16857), .SI(test_si100), .SE(test_se), .CLK(CK), 
        .Q(g8271), .QN() );
  SDFFX1 DFF_1622_Q_reg ( .D(g16866), .SI(g8271), .SE(test_se), .CLK(CK), .Q(
        g3083), .QN() );
  SDFFX1 DFF_1623_Q_reg ( .D(n4261), .SI(g3083), .SE(test_se), .CLK(CK), .Q(
        g8267), .QN() );
  SDFFX1 DFF_1624_Q_reg ( .D(N995), .SI(g8267), .SE(test_se), .CLK(CK), .Q(
        n4577), .QN() );
  SDFFX1 DFF_1625_Q_reg ( .D(g16845), .SI(n4577), .SE(test_se), .CLK(CK), .Q(
        g8266), .QN(DFF_1625_n1) );
  SDFFX1 DFF_1626_Q_reg ( .D(g16854), .SI(g8266), .SE(test_se), .CLK(CK), .Q(
        g8265), .QN(DFF_1626_n1) );
  SDFFX1 DFF_1627_Q_reg ( .D(g16861), .SI(g8265), .SE(test_se), .CLK(CK), .Q(
        g8264), .QN() );
  SDFFX1 DFF_1628_Q_reg ( .D(g16880), .SI(g8264), .SE(test_se), .CLK(CK), .Q(
        g8262), .QN(DFF_1628_n1) );
  SDFFX1 DFF_1629_Q_reg ( .D(g18755), .SI(g8262), .SE(test_se), .CLK(CK), .Q(
        g8263), .QN() );
  SDFFX1 DFF_1630_Q_reg ( .D(g18804), .SI(g8263), .SE(test_se), .CLK(CK), .Q(
        g8260), .QN() );
  SDFFX1 DFF_1631_Q_reg ( .D(g18837), .SI(g8260), .SE(test_se), .CLK(CK), .Q(
        g8261), .QN() );
  SDFFX1 DFF_1632_Q_reg ( .D(g18868), .SI(g8261), .SE(test_se), .CLK(CK), .Q(
        g8259), .QN() );
  SDFFX1 DFF_1633_Q_reg ( .D(g18907), .SI(g8259), .SE(test_se), .CLK(CK), .Q(
        g2990), .QN() );
  SDFFX1 DFF_1634_Q_reg ( .D(N690), .SI(g2990), .SE(test_se), .CLK(CK), .Q(
        n4578), .QN() );
  SDFFX1 DFF_1635_Q_reg ( .D(n4260), .SI(n4578), .SE(test_se), .CLK(CK), .Q(
        g8258), .QN() );
  SDFFX1 DFF_454_Q_reg ( .D(n4598), .SI(n8040), .SE(test_se), .CLK(CK), .Q(
        g6677), .QN(n4309) );
  SDFFX1 DFF_804_Q_reg ( .D(n4598), .SI(test_si49), .SE(test_se), .CLK(CK), 
        .Q(g6979), .QN(n4308) );
  SDFFX1 DFF_1154_Q_reg ( .D(n4598), .SI(n7960), .SE(test_se), .CLK(CK), .Q(
        g7229), .QN(n4307) );
  SDFFX1 DFF_1504_Q_reg ( .D(n4597), .SI(n7918), .SE(test_se), .CLK(CK), .Q(
        g7425), .QN(n4306) );
  SDFFX1 DFF_1300_Q_reg ( .D(n4610), .SI(g2351), .SE(test_se), .CLK(CK), .Q(
        g2480), .QN(n4524) );
  SDFFX1 DFF_950_Q_reg ( .D(n4622), .SI(g1657), .SE(test_se), .CLK(CK), .Q(
        g1786), .QN(n4525) );
  SDFFX1 DFF_951_Q_reg ( .D(n4620), .SI(g1786), .SE(test_se), .CLK(CK), .Q(
        g1782), .QN(n4511) );
  SDFFX1 DFF_1301_Q_reg ( .D(n4608), .SI(g2480), .SE(test_se), .CLK(CK), .Q(
        g2476), .QN(n4509) );
  SDFFX1 DFF_250_Q_reg ( .D(n4643), .SI(g276), .SE(test_se), .CLK(CK), .Q(
        g6447), .QN(n4499) );
  SDFFX1 DFF_249_Q_reg ( .D(n4650), .SI(g181), .SE(test_se), .CLK(CK), .Q(g276), .QN(n4520) );
  NAND3X1 U3788 ( .IN1(n2773), .IN2(n2774), .IN3(n2775), .QN(n2718) );
  NAND3X1 U3789 ( .IN1(n2734), .IN2(n2735), .IN3(n2736), .QN(n2670) );
  NAND3X1 U3790 ( .IN1(n2749), .IN2(n2750), .IN3(n2751), .QN(n2685) );
  INVX0 U3791 ( .IN(n2513), .QN(n2077) );
  INVX0 U3792 ( .IN(n2539), .QN(n1975) );
  NAND2X0 U3793 ( .IN1(n1791), .IN2(n1787), .QN(n2720) );
  INVX0 U3794 ( .IN(n2591), .QN(n1769) );
  AND2X1 U3795 ( .IN1(n2720), .IN2(n2569), .Q(n4507) );
  INVX0 U3796 ( .IN(n2823), .QN(n2099) );
  INVX0 U3797 ( .IN(n2498), .QN(n2079) );
  OA222X1 U3798 ( .IN1(n4524), .IN2(g2394), .IN3(n4509), .IN4(g2395), .IN5(
        n4516), .IN6(g2393), .Q(n2787) );
  NAND2X0 U3799 ( .IN1(n2787), .IN2(n4116), .QN(n2823) );
  INVX0 U3800 ( .IN(n2778), .QN(n2095) );
  NAND2X0 U3801 ( .IN1(n3683), .IN2(g2147), .QN(n3425) );
  NAND2X0 U3802 ( .IN1(n3887), .IN2(test_so78), .QN(n3684) );
  NAND2X0 U3803 ( .IN1(n2099), .IN2(n2095), .QN(n2672) );
  AOI222X1 U3804 ( .IN1(g2345), .IN2(n4587), .IN3(g2348), .IN4(n4679), .IN5(
        g2342), .IN6(g6837), .QN(n2499) );
  INVX0 U3805 ( .IN(n4517), .QN(n2725) );
  INVX0 U3806 ( .IN(n2833), .QN(n1997) );
  INVX0 U3807 ( .IN(n2525), .QN(n1977) );
  OA222X1 U3808 ( .IN1(n4525), .IN2(g1700), .IN3(n4511), .IN4(g1701), .IN5(
        n4518), .IN6(g1699), .Q(n2606) );
  NAND2X0 U3809 ( .IN1(n2606), .IN2(n4117), .QN(n2833) );
  INVX0 U3810 ( .IN(n2597), .QN(n1993) );
  NAND2X0 U3811 ( .IN1(n3686), .IN2(g1453), .QN(n3428) );
  NAND2X0 U3812 ( .IN1(n3890), .IN2(g1462), .QN(n3687) );
  NAND2X0 U3813 ( .IN1(n1997), .IN2(n1993), .QN(n2687) );
  INVX0 U3814 ( .IN(n4519), .QN(n2741) );
  INVX0 U3815 ( .IN(n2813), .QN(n1791) );
  INVX0 U3816 ( .IN(n2577), .QN(n1771) );
  OA222X1 U3817 ( .IN1(n4676), .IN2(g319), .IN3(n4506), .IN4(g320), .IN5(n4520), .IN6(g318), .Q(n2647) );
  NAND2X0 U3818 ( .IN1(n2647), .IN2(n4119), .QN(n2813) );
  NAND2X0 U3819 ( .IN1(n3692), .IN2(test_so15), .QN(n3434) );
  NAND2X0 U3820 ( .IN1(n3896), .IN2(g88), .QN(n3693) );
  NBUFFX2 U3821 ( .IN(n2720), .Q(n4498) );
  NAND2X0 U3822 ( .IN1(g186), .IN2(g138), .QN(n4497) );
  NAND2X0 U3823 ( .IN1(test_so13), .IN2(g6313), .QN(n4495) );
  NAND2X0 U3824 ( .IN1(g192), .IN2(n4694), .QN(n4496) );
  INVX0 U3825 ( .IN(n4507), .QN(n2771) );
  NBUFFX2 U3826 ( .IN(n4499), .Q(n4676) );
  INVX0 U3827 ( .IN(g2241), .QN(n4680) );
  INVX0 U3828 ( .IN(n4680), .QN(n4679) );
  INVX0 U3829 ( .IN(g1547), .QN(n4685) );
  INVX0 U3830 ( .IN(n4685), .QN(n4684) );
  INVX0 U3831 ( .IN(g165), .QN(n4695) );
  INVX0 U3832 ( .IN(n4695), .QN(n4694) );
  INVX0 U3833 ( .IN(n2720), .QN(n1785) );
  INVX0 U3834 ( .IN(n2638), .QN(n1787) );
  INVX0 U3835 ( .IN(n4324), .QN(g6837) );
  INVX0 U3836 ( .IN(n4317), .QN(g6573) );
  INVX0 U3837 ( .IN(n4318), .QN(g6231) );
  NAND3X0 U3838 ( .IN1(n4495), .IN2(n4496), .IN3(n4497), .QN(n2591) );
  AND2X1 U3839 ( .IN1(n2099), .IN2(n2095), .Q(n4508) );
  AND2X1 U3840 ( .IN1(n1997), .IN2(n1993), .Q(n4510) );
  NAND2X0 U3841 ( .IN1(g2261), .IN2(g2214), .QN(n4502) );
  NAND2X0 U3842 ( .IN1(g1567), .IN2(g1520), .QN(n4505) );
  NAND2X0 U3843 ( .IN1(test_so76), .IN2(g7084), .QN(n4500) );
  NAND2X0 U3844 ( .IN1(g2267), .IN2(n4679), .QN(n4501) );
  NAND3X0 U3845 ( .IN1(n4500), .IN2(n4501), .IN3(n4502), .QN(n2513) );
  NAND2X0 U3846 ( .IN1(g1570), .IN2(g6782), .QN(n4503) );
  NAND2X0 U3847 ( .IN1(g1573), .IN2(n4684), .QN(n4504) );
  NAND3X0 U3848 ( .IN1(n4503), .IN2(n4504), .IN3(n4505), .QN(n2539) );
  LSDNX1 U3849 ( .D(n1769), .Q(n4513) );
  NAND2X0 U3850 ( .IN1(n4694), .IN2(n4652), .QN(n3897) );
  AND2X1 U3851 ( .IN1(n2672), .IN2(n2490), .Q(n4517) );
  AND2X1 U3852 ( .IN1(n2687), .IN2(n2517), .Q(n4519) );
  OR2X1 U3853 ( .IN1(n3424), .IN2(g2138), .Q(n3423) );
  OR2X1 U3854 ( .IN1(n3427), .IN2(g1444), .Q(n3426) );
  OR2X1 U3855 ( .IN1(n3433), .IN2(g70), .Q(n3432) );
  LSDNX1 U3856 ( .D(n4508), .Q(n4529) );
  LSDNX1 U3857 ( .D(n4510), .Q(n4530) );
  NBUFFX2 U3858 ( .IN(n2505), .Q(n4651) );
  NBUFFX2 U3859 ( .IN(n2505), .Q(n4652) );
  LSDNX1 U3860 ( .D(n3425), .Q(n4522) );
  LSDNX1 U3861 ( .D(n3428), .Q(n4523) );
  LSDNX1 U3862 ( .D(n3434), .Q(n4521) );
  NAND2X1 U3863 ( .IN1(n3171), .IN2(g61), .QN(n2991) );
  NAND2X1 U3864 ( .IN1(n3159), .IN2(g2129), .QN(n2982) );
  NAND2X1 U3865 ( .IN1(n3163), .IN2(g1435), .QN(n2985) );
  INVX0 U3866 ( .IN(n2292), .QN(n1568) );
  NOR2X0 U3867 ( .IN1(g2896), .IN2(g2892), .QN(n4223) );
  NAND2X0 U3868 ( .IN1(n3893), .IN2(g776), .QN(n3690) );
  NAND2X0 U3869 ( .IN1(n3689), .IN2(g767), .QN(n3431) );
  NAND2X0 U3870 ( .IN1(n3430), .IN2(g758), .QN(n3168) );
  NBUFFX2 U3871 ( .IN(g545), .Q(n4638) );
  NAND2X0 U3872 ( .IN1(n3424), .IN2(g2138), .QN(n3160) );
  NAND2X0 U3873 ( .IN1(n3427), .IN2(g1444), .QN(n3164) );
  NAND2X0 U3874 ( .IN1(n3433), .IN2(g70), .QN(n3172) );
  OR2X1 U3875 ( .IN1(n3430), .IN2(g758), .Q(n3429) );
  OR2X1 U3876 ( .IN1(n3689), .IN2(g767), .Q(n3688) );
  OR2X1 U3877 ( .IN1(n3893), .IN2(g776), .Q(n3892) );
  OR2X1 U3878 ( .IN1(n3683), .IN2(g2147), .Q(n3682) );
  OR2X1 U3879 ( .IN1(n3686), .IN2(g1453), .Q(n3685) );
  OR2X1 U3880 ( .IN1(n3692), .IN2(test_so15), .Q(n3691) );
  LSDNX1 U3881 ( .D(g1231), .Q(g6750) );
  AO222X1 U3882 ( .IN1(test_so77), .IN2(n4587), .IN3(g2330), .IN4(n4679), 
        .IN5(g2324), .IN6(g6837), .Q(n2503) );
  AO222X1 U3883 ( .IN1(g1633), .IN2(n4589), .IN3(g1636), .IN4(n4684), .IN5(
        g1630), .IN6(g6573), .Q(n2530) );
  AO222X1 U3884 ( .IN1(g252), .IN2(n4593), .IN3(test_so14), .IN4(n4694), .IN5(
        g249), .IN6(g6231), .Q(n2582) );
  AO222X1 U3885 ( .IN1(g2318), .IN2(n4587), .IN3(g2321), .IN4(n4679), .IN5(
        g2315), .IN6(g6837), .Q(n2708) );
  AO222X1 U3886 ( .IN1(g1624), .IN2(n4589), .IN3(g1627), .IN4(n4684), .IN5(
        test_so55), .IN6(g6573), .Q(n2727) );
  AO222X1 U3887 ( .IN1(g243), .IN2(n4593), .IN3(g246), .IN4(n4694), .IN5(g240), 
        .IN6(g6231), .Q(n2759) );
  LSDNX1 U3888 ( .D(n3687), .Q(n4527) );
  LSDNX1 U3889 ( .D(n3693), .Q(n4528) );
  LSDNX1 U3890 ( .D(n3684), .Q(n4526) );
  NORI3X1 U3891 ( .IN1(g1943), .IN2(g1939), .IN3(n1818), .QN(n2313) );
  NAND2X1 U3892 ( .IN1(n3167), .IN2(test_so36), .QN(n2988) );
  NAND2X0 U3893 ( .IN1(test_so31), .IN2(n4651), .QN(n3894) );
  NAND2X0 U3894 ( .IN1(n4679), .IN2(n4652), .QN(n3888) );
  NAND2X0 U3895 ( .IN1(n4684), .IN2(n4652), .QN(n3891) );
  INVX0 U3896 ( .IN(n2454), .QN(n1583) );
  INVX0 U3897 ( .IN(n2364), .QN(n1570) );
  INVX0 U3898 ( .IN(n2220), .QN(n1566) );
  INVX0 U3899 ( .IN(n2363), .QN(n2136) );
  INVX0 U3900 ( .IN(n2219), .QN(n1932) );
  LSDNENX1 U3901 ( .D(n2302), .ENB(n2289), .Q(n2303) );
  LSDNENX1 U3902 ( .D(n2313), .ENB(n2289), .Q(n2275) );
  INVX0 U3903 ( .IN(n2291), .QN(n2034) );
  NAND2X0 U3904 ( .IN1(n2472), .IN2(n2473), .QN(n2451) );
  NAND2X0 U3905 ( .IN1(n2394), .IN2(n2395), .QN(n2388) );
  NAND2X0 U3906 ( .IN1(n2250), .IN2(n2251), .QN(n2244) );
  NAND2X0 U3907 ( .IN1(n2322), .IN2(n2323), .QN(n2316) );
  INVX0 U3908 ( .IN(n2439), .QN(n1584) );
  INVX0 U3909 ( .IN(n2384), .QN(n2154) );
  INVX0 U3910 ( .IN(n2312), .QN(n2052) );
  INVX0 U3911 ( .IN(n2240), .QN(n1950) );
  INVX0 U3912 ( .IN(n2444), .QN(n1849) );
  INVX0 U3913 ( .IN(n2373), .QN(n2155) );
  INVX0 U3914 ( .IN(n2301), .QN(n2053) );
  INVX0 U3915 ( .IN(n2229), .QN(n1951) );
  INVX0 U3916 ( .IN(n2448), .QN(n1850) );
  INVX0 U3917 ( .IN(n2442), .QN(n1847) );
  INVX0 U3918 ( .IN(n2377), .QN(n2152) );
  INVX0 U3919 ( .IN(n2305), .QN(n2050) );
  INVX0 U3920 ( .IN(n2233), .QN(n1948) );
  INVX0 U3921 ( .IN(n2471), .QN(n1855) );
  INVX0 U3922 ( .IN(n2382), .QN(n2160) );
  INVX0 U3923 ( .IN(n2310), .QN(n2058) );
  INVX0 U3924 ( .IN(n2238), .QN(n1956) );
  INVX0 U3925 ( .IN(n2431), .QN(n1851) );
  INVX0 U3926 ( .IN(n2352), .QN(n2156) );
  INVX0 U3927 ( .IN(n2280), .QN(n2054) );
  INVX0 U3928 ( .IN(n2208), .QN(n1952) );
  INVX0 U3929 ( .IN(n2464), .QN(n1854) );
  INVX0 U3930 ( .IN(n2368), .QN(n2159) );
  INVX0 U3931 ( .IN(n2296), .QN(n2057) );
  INVX0 U3932 ( .IN(n2224), .QN(n1955) );
  INVX0 U3933 ( .IN(n2360), .QN(n1569) );
  INVX0 U3934 ( .IN(n2216), .QN(n1565) );
  NAND2X0 U3935 ( .IN1(g2993), .IN2(n4597), .QN(n3859) );
  NAND2X0 U3936 ( .IN1(g3006), .IN2(n4130), .QN(n4066) );
  NAND2X0 U3937 ( .IN1(n2313), .IN2(g1880), .QN(n2288) );
  NAND2X0 U3938 ( .IN1(n2426), .IN2(n2427), .QN(n4265) );
  OR2X1 U3939 ( .IN1(n4065), .IN2(g3013), .Q(n4064) );
  OR2X1 U3940 ( .IN1(n3167), .IN2(test_so36), .Q(n3166) );
  OR2X1 U3941 ( .IN1(n3159), .IN2(g2129), .Q(n3158) );
  OR2X1 U3942 ( .IN1(n3163), .IN2(g1435), .Q(n3162) );
  OR2X1 U3943 ( .IN1(n3171), .IN2(g61), .Q(n3170) );
  AOI21X1 U3944 ( .IN1(g2574), .IN2(DFF_1449_n1), .IN3(n2960), .QN(g30072) );
  OR2X1 U3945 ( .IN1(n4130), .IN2(g3006), .Q(n4128) );
  OR2X1 U3946 ( .IN1(n3887), .IN2(test_so78), .Q(n3886) );
  OR2X1 U3947 ( .IN1(n3890), .IN2(g1462), .Q(n3889) );
  OR2X1 U3948 ( .IN1(n3896), .IN2(g88), .Q(n3895) );
  XOR3X1 U3949 ( .IN1(n2414), .IN2(n4531), .IN3(n2416), .Q(n2407) );
  XOR2X1 U3950 ( .IN1(n2417), .IN2(n2418), .Q(n4531) );
  XNOR3X1 U3951 ( .IN1(n2337), .IN2(n4532), .IN3(n2339), .Q(n2336) );
  XOR2X1 U3952 ( .IN1(n2340), .IN2(n2341), .Q(n4532) );
  XNOR3X1 U3953 ( .IN1(n2265), .IN2(n4533), .IN3(n2267), .Q(n2264) );
  XOR2X1 U3954 ( .IN1(n2268), .IN2(n2269), .Q(n4533) );
  XNOR3X1 U3955 ( .IN1(n2193), .IN2(n4534), .IN3(n2195), .Q(n2192) );
  XOR2X1 U3956 ( .IN1(n2196), .IN2(n2197), .Q(n4534) );
  NOR2X2 U3957 ( .IN1(n2293), .IN2(n2034), .QN(n2289) );
  NOR2X0 U3958 ( .IN1(n4535), .IN2(n2777), .QN(n2592) );
  XNOR2X1 U3959 ( .IN1(n2778), .IN2(n2779), .Q(n4535) );
  NOR2X0 U3960 ( .IN1(n4536), .IN2(n2596), .QN(n2593) );
  XNOR2X1 U3961 ( .IN1(n2597), .IN2(n2598), .Q(n4536) );
  NOR2X0 U3962 ( .IN1(n4537), .IN2(n2637), .QN(n2615) );
  XNOR2X1 U3963 ( .IN1(n2638), .IN2(n2639), .Q(n4537) );
  NOR2X0 U3964 ( .IN1(n4538), .IN2(n2777), .QN(n2796) );
  XNOR2X1 U3965 ( .IN1(n2821), .IN2(n2787), .Q(n4538) );
  NOR2X0 U3966 ( .IN1(n4539), .IN2(n2596), .QN(n2797) );
  XNOR2X1 U3967 ( .IN1(n2831), .IN2(n2606), .Q(n4539) );
  NOR2X0 U3968 ( .IN1(n4540), .IN2(n2637), .QN(n2799) );
  XNOR2X1 U3969 ( .IN1(n2811), .IN2(n2647), .Q(n4540) );
  INVX0 U3970 ( .IN(n2385), .QN(n4552) );
  INVX0 U3971 ( .IN(n2241), .QN(n4551) );
  OR2X1 U3972 ( .IN1(n4541), .IN2(n4542), .Q(n2445) );
  OA221X1 U3973 ( .IN1(n4359), .IN2(g736), .IN3(n4295), .IN4(g734), .IN5(n2450), .Q(n4542) );
  OR2X1 U3974 ( .IN1(n4543), .IN2(n4544), .Q(n2374) );
  OA221X1 U3975 ( .IN1(n4356), .IN2(g2810), .IN3(n4292), .IN4(g2808), .IN5(
        n2387), .Q(n4544) );
  OR2X1 U3976 ( .IN1(n4545), .IN2(n4546), .Q(n2302) );
  OA221X1 U3977 ( .IN1(n4357), .IN2(g2116), .IN3(n4293), .IN4(g2114), .IN5(
        n2315), .Q(n4546) );
  OR2X1 U3978 ( .IN1(n4548), .IN2(n4547), .Q(n2230) );
  OA221X1 U3979 ( .IN1(n4358), .IN2(g1422), .IN3(n4294), .IN4(g1420), .IN5(
        n2243), .Q(n4547) );
  OAI21X1 U3980 ( .IN1(n4548), .IN2(n4549), .IN3(n4550), .QN(n3156) );
  AO221X1 U3981 ( .IN1(n4371), .IN2(n4361), .IN3(g21851), .IN4(g6750), .IN5(
        g1186), .Q(n4550) );
  NAND2X1 U3982 ( .IN1(n4065), .IN2(g3013), .QN(n3742) );
  LSDNX1 U3983 ( .D(g1925), .Q(g7052) );
  LSDNX1 U3984 ( .D(g2619), .Q(g7302) );
  LSDNX1 U3985 ( .D(g2480), .Q(n4608) );
  LSDNX1 U3986 ( .D(g1786), .Q(n4620) );
  LSDNX1 U3987 ( .D(g6447), .Q(n4641) );
  LSDNX1 U3988 ( .D(g545), .Q(g6485) );
  LSDNX1 U3989 ( .D(g2351), .Q(n4610) );
  LSDNX1 U3990 ( .D(g1657), .Q(n4622) );
  LSDNX1 U3991 ( .D(g276), .Q(n4643) );
  LSDNX1 U3992 ( .D(g2476), .Q(n4606) );
  LSDNX1 U3993 ( .D(g1782), .Q(n4618) );
  LSDNX1 U3994 ( .D(g401), .Q(n4640) );
  LSDNX1 U3995 ( .D(g3080), .Q(n4598) );
  NAND2X0 U3996 ( .IN1(n4551), .IN2(n2217), .QN(n2203) );
  NAND2X0 U3997 ( .IN1(n4552), .IN2(n2361), .QN(n2347) );
  NOR4X1 U3998 ( .IN1(g21851), .IN2(n2480), .IN3(g563), .IN4(g559), .QN(n2478)
         );
  NOR2X2 U3999 ( .IN1(n2455), .IN2(n1832), .QN(n2446) );
  INVX0 U4000 ( .IN(n4754), .QN(n4736) );
  INVX0 U4001 ( .IN(n4753), .QN(n4737) );
  INVX0 U4002 ( .IN(n4753), .QN(n4734) );
  INVX0 U4003 ( .IN(n4753), .QN(n4735) );
  NOR2X0 U4004 ( .IN1(n1689), .IN2(n2661), .QN(n2659) );
  NOR2X0 U4005 ( .IN1(n1632), .IN2(n2675), .QN(n2673) );
  NOR2X0 U4006 ( .IN1(n1651), .IN2(n2690), .QN(n2688) );
  NOR2X0 U4007 ( .IN1(n1670), .IN2(n2704), .QN(n2702) );
  NOR2X0 U4008 ( .IN1(n2722), .IN2(n2672), .QN(n2668) );
  NOR2X0 U4009 ( .IN1(n2738), .IN2(n2687), .QN(n2683) );
  NOR2X0 U4010 ( .IN1(n2768), .IN2(n4498), .QN(n2716) );
  NOR2X0 U4011 ( .IN1(n2753), .IN2(n2754), .QN(n2698) );
  INVX0 U4012 ( .IN(n4763), .QN(n4753) );
  INVX0 U4013 ( .IN(n4762), .QN(n4754) );
  NOR2X0 U4014 ( .IN1(n2722), .IN2(n4529), .QN(n2662) );
  NOR2X0 U4015 ( .IN1(n2738), .IN2(n4530), .QN(n2676) );
  NOR2X0 U4016 ( .IN1(n2753), .IN2(n1889), .QN(n2691) );
  NOR2X0 U4017 ( .IN1(n2768), .IN2(n1785), .QN(n2705) );
  INVX0 U4018 ( .IN(n2661), .QN(n1688) );
  INVX0 U4019 ( .IN(n2675), .QN(n1631) );
  INVX0 U4020 ( .IN(n2690), .QN(n1650) );
  INVX0 U4021 ( .IN(n2704), .QN(n1669) );
  INVX0 U4022 ( .IN(n2754), .QN(n1889) );
  INVX0 U4023 ( .IN(n2722), .QN(n1689) );
  INVX0 U4024 ( .IN(n2738), .QN(n1632) );
  INVX0 U4025 ( .IN(n2753), .QN(n1651) );
  INVX0 U4026 ( .IN(n2768), .QN(n1670) );
  INVX0 U4027 ( .IN(n4700), .QN(n4731) );
  INVX0 U4028 ( .IN(n4768), .QN(n4741) );
  INVX0 U4029 ( .IN(n4769), .QN(n4740) );
  INVX0 U4030 ( .IN(n4769), .QN(n4739) );
  INVX0 U4031 ( .IN(n4768), .QN(n4742) );
  INVX0 U4032 ( .IN(n4767), .QN(n4744) );
  INVX0 U4033 ( .IN(n4766), .QN(n4746) );
  INVX0 U4034 ( .IN(n4766), .QN(n4745) );
  INVX0 U4035 ( .IN(n4765), .QN(n4749) );
  INVX0 U4036 ( .IN(n4765), .QN(n4748) );
  INVX0 U4037 ( .IN(n4766), .QN(n4747) );
  INVX0 U4038 ( .IN(n4764), .QN(n4751) );
  INVX0 U4039 ( .IN(n4764), .QN(n4750) );
  INVX0 U4040 ( .IN(n4763), .QN(n4752) );
  INVX0 U4041 ( .IN(n4762), .QN(n4755) );
  INVX0 U4042 ( .IN(n4761), .QN(n4756) );
  INVX0 U4043 ( .IN(n4761), .QN(n4757) );
  INVX0 U4044 ( .IN(n4760), .QN(n4758) );
  INVX0 U4045 ( .IN(n4721), .QN(n4706) );
  INVX0 U4046 ( .IN(n4721), .QN(n4707) );
  INVX0 U4047 ( .IN(n4722), .QN(n4705) );
  INVX0 U4048 ( .IN(n4722), .QN(n4704) );
  INVX0 U4049 ( .IN(n4723), .QN(n4703) );
  INVX0 U4050 ( .IN(n4723), .QN(n4702) );
  INVX0 U4051 ( .IN(n4720), .QN(n4708) );
  INVX0 U4052 ( .IN(n4718), .QN(n4712) );
  INVX0 U4053 ( .IN(n4720), .QN(n4709) );
  INVX0 U4054 ( .IN(n4717), .QN(n4715) );
  INVX0 U4055 ( .IN(n4717), .QN(n4714) );
  INVX0 U4056 ( .IN(n4718), .QN(n4713) );
  INVX0 U4057 ( .IN(n4719), .QN(n4711) );
  INVX0 U4058 ( .IN(n4719), .QN(n4710) );
  INVX0 U4059 ( .IN(n4351), .QN(n4716) );
  INVX0 U4060 ( .IN(n4760), .QN(n4759) );
  INVX0 U4061 ( .IN(n3161), .QN(n1605) );
  INVX0 U4062 ( .IN(n3165), .QN(n1604) );
  INVX0 U4063 ( .IN(n3169), .QN(n1603) );
  INVX0 U4064 ( .IN(n3157), .QN(n1606) );
  XOR3X1 U4065 ( .IN1(n2409), .IN2(n2410), .IN3(n2411), .Q(n2408) );
  XOR2X1 U4066 ( .IN1(n2412), .IN2(n2413), .Q(n2410) );
  AO221X1 U4067 ( .IN1(n2659), .IN2(n2081), .IN3(n2733), .IN4(n2661), .IN5(
        n2662), .Q(n2711) );
  XOR2X1 U4068 ( .IN1(n2670), .IN2(n2080), .Q(n2733) );
  AO221X1 U4069 ( .IN1(n2673), .IN2(n1979), .IN3(n2748), .IN4(n2675), .IN5(
        n2676), .Q(n2730) );
  XOR2X1 U4070 ( .IN1(n2685), .IN2(n1978), .Q(n2748) );
  AO221X1 U4071 ( .IN1(n2702), .IN2(n1773), .IN3(n2772), .IN4(n2704), .IN5(
        n2705), .Q(n2762) );
  XOR2X1 U4072 ( .IN1(n2718), .IN2(n1772), .Q(n2772) );
  XOR2X1 U4073 ( .IN1(n4508), .IN2(n2079), .Q(n2710) );
  XOR2X1 U4074 ( .IN1(n4510), .IN2(n1977), .Q(n2729) );
  XOR2X1 U4075 ( .IN1(n1785), .IN2(n1771), .Q(n2761) );
  XOR2X1 U4076 ( .IN1(n4508), .IN2(n2077), .Q(n2724) );
  XOR2X1 U4077 ( .IN1(n4510), .IN2(n1975), .Q(n2740) );
  XOR2X1 U4078 ( .IN1(n1785), .IN2(n1769), .Q(n2770) );
  XOR3X1 U4079 ( .IN1(n2342), .IN2(n2343), .IN3(n2344), .Q(n2335) );
  XNOR2X1 U4080 ( .IN1(n2345), .IN2(n2346), .Q(n2343) );
  XOR3X1 U4081 ( .IN1(n2270), .IN2(n2271), .IN3(n2272), .Q(n2263) );
  XNOR2X1 U4082 ( .IN1(n2273), .IN2(n2274), .Q(n2271) );
  NOR2X0 U4083 ( .IN1(n1766), .IN2(n4553), .QN(n4074) );
  NOR2X0 U4084 ( .IN1(n1765), .IN2(n4553), .QN(n4075) );
  NOR2X0 U4085 ( .IN1(n1764), .IN2(n4553), .QN(n4076) );
  NOR2X0 U4086 ( .IN1(n1763), .IN2(n4553), .QN(n4079) );
  NOR2X0 U4087 ( .IN1(n1762), .IN2(n4553), .QN(n4080) );
  NOR2X0 U4088 ( .IN1(n1761), .IN2(n4553), .QN(n4085) );
  NOR2X0 U4089 ( .IN1(n1760), .IN2(n4553), .QN(n4086) );
  NOR2X0 U4090 ( .IN1(n1759), .IN2(n4553), .QN(n4091) );
  NAND3X0 U4091 ( .IN1(n1854), .IN2(n1851), .IN3(n1855), .QN(n2474) );
  NAND3X0 U4092 ( .IN1(n2159), .IN2(n2156), .IN3(n2160), .QN(n2396) );
  NAND3X0 U4093 ( .IN1(n2057), .IN2(n2054), .IN3(n2058), .QN(n2324) );
  NAND3X0 U4094 ( .IN1(n1955), .IN2(n1952), .IN3(n1956), .QN(n2252) );
  XOR3X1 U4095 ( .IN1(n2198), .IN2(n2199), .IN3(n2200), .Q(n2191) );
  XNOR2X1 U4096 ( .IN1(n2201), .IN2(n2202), .Q(n2199) );
  INVX0 U4097 ( .IN(n3740), .QN(n1581) );
  INVX0 U4098 ( .IN(n3503), .QN(n2122) );
  INVX0 U4099 ( .IN(n3504), .QN(n2123) );
  INVX0 U4100 ( .IN(n3508), .QN(n2121) );
  INVX0 U4101 ( .IN(n3507), .QN(n2020) );
  INVX0 U4102 ( .IN(n3514), .QN(n2021) );
  INVX0 U4103 ( .IN(n3525), .QN(n2019) );
  INVX0 U4104 ( .IN(n3517), .QN(n1918) );
  INVX0 U4105 ( .IN(n3531), .QN(n1919) );
  INVX0 U4106 ( .IN(n3551), .QN(n1917) );
  INVX0 U4107 ( .IN(n3534), .QN(n1814) );
  INVX0 U4108 ( .IN(n3557), .QN(n1815) );
  INVX0 U4109 ( .IN(n3586), .QN(n1813) );
  OA21X1 U4110 ( .IN1(n4517), .IN2(n2894), .IN3(n2892), .Q(n2661) );
  OA21X1 U4111 ( .IN1(n4529), .IN2(n2489), .IN3(n2893), .Q(n2894) );
  OA21X1 U4112 ( .IN1(n4519), .IN2(n2912), .IN3(n2910), .Q(n2675) );
  OA21X1 U4113 ( .IN1(n4530), .IN2(n2516), .IN3(n2911), .Q(n2912) );
  OA21X1 U4114 ( .IN1(n1890), .IN2(n2930), .IN3(n2928), .Q(n2690) );
  INVX0 U4115 ( .IN(n2757), .QN(n1890) );
  OA21X1 U4116 ( .IN1(n1889), .IN2(n2542), .IN3(n2929), .Q(n2930) );
  OA21X1 U4117 ( .IN1(n4507), .IN2(n2947), .IN3(n2945), .Q(n2704) );
  OA21X1 U4118 ( .IN1(n1785), .IN2(n2568), .IN3(n2946), .Q(n2947) );
  NAND2X0 U4119 ( .IN1(n1895), .IN2(n1891), .QN(n2754) );
  NAND2X0 U4120 ( .IN1(n2754), .IN2(n2543), .QN(n2757) );
  NOR2X0 U4121 ( .IN1(n4654), .IN2(n1845), .QN(n2433) );
  NOR2X0 U4122 ( .IN1(n4660), .IN2(n2150), .QN(n2354) );
  NOR2X0 U4123 ( .IN1(n4658), .IN2(n2048), .QN(n2282) );
  NOR2X0 U4124 ( .IN1(n4656), .IN2(n1946), .QN(n2210) );
  NOR2X0 U4125 ( .IN1(n2829), .IN2(n2899), .QN(n2790) );
  NOR2X0 U4126 ( .IN1(n2839), .IN2(n2917), .QN(n2609) );
  NOR2X0 U4127 ( .IN1(n2809), .IN2(n2935), .QN(n2630) );
  NOR2X0 U4128 ( .IN1(n2819), .IN2(n2952), .QN(n2650) );
  NOR2X0 U4129 ( .IN1(n4653), .IN2(n1845), .QN(n2438) );
  NOR2X0 U4130 ( .IN1(n4659), .IN2(n2150), .QN(n2359) );
  NOR2X0 U4131 ( .IN1(n4657), .IN2(n2048), .QN(n2287) );
  NOR2X0 U4132 ( .IN1(n4655), .IN2(n1946), .QN(n2215) );
  NAND3X0 U4133 ( .IN1(n2891), .IN2(n2725), .IN3(n2892), .QN(n2722) );
  NAND2X0 U4134 ( .IN1(n2489), .IN2(n2893), .QN(n2891) );
  NAND3X0 U4135 ( .IN1(n2909), .IN2(n2741), .IN3(n2910), .QN(n2738) );
  NAND2X0 U4136 ( .IN1(n2516), .IN2(n2911), .QN(n2909) );
  NAND3X0 U4137 ( .IN1(n2927), .IN2(n2757), .IN3(n2928), .QN(n2753) );
  NAND2X0 U4138 ( .IN1(n2542), .IN2(n2929), .QN(n2927) );
  NAND3X0 U4139 ( .IN1(n2944), .IN2(n2771), .IN3(n2945), .QN(n2768) );
  NAND2X0 U4140 ( .IN1(n2568), .IN2(n2946), .QN(n2944) );
  INVX0 U4141 ( .IN(n4774), .QN(n4763) );
  INVX0 U4142 ( .IN(n4774), .QN(n4762) );
  XOR2X1 U4143 ( .IN1(n1889), .IN2(n1876), .Q(n2745) );
  XOR2X1 U4144 ( .IN1(n1889), .IN2(n1874), .Q(n2756) );
  INVX0 U4145 ( .IN(n2899), .QN(n1687) );
  INVX0 U4146 ( .IN(n2917), .QN(n1630) );
  INVX0 U4147 ( .IN(n2935), .QN(n1649) );
  INVX0 U4148 ( .IN(n2952), .QN(n1668) );
  NAND2X0 U4149 ( .IN1(n2789), .IN2(n2794), .QN(n2829) );
  NAND2X0 U4150 ( .IN1(n2608), .IN2(n2613), .QN(n2839) );
  NAND2X0 U4151 ( .IN1(n2629), .IN2(n2634), .QN(n2809) );
  NAND2X0 U4152 ( .IN1(n2649), .IN2(n2654), .QN(n2819) );
  AO21X1 U4153 ( .IN1(n2119), .IN2(n3281), .IN3(n2117), .Q(n3280) );
  NAND2X0 U4154 ( .IN1(n2118), .IN2(n2129), .QN(n3281) );
  INVX0 U4155 ( .IN(n3282), .QN(n2117) );
  NBUFFX2 U4156 ( .IN(n4364), .Q(n4671) );
  NBUFFX2 U4157 ( .IN(n4363), .Q(n4673) );
  NBUFFX2 U4158 ( .IN(n4381), .Q(n4669) );
  NBUFFX2 U4159 ( .IN(n4524), .Q(n4664) );
  NBUFFX2 U4160 ( .IN(n4525), .Q(n4667) );
  NBUFFX2 U4161 ( .IN(n4364), .Q(n4672) );
  NBUFFX2 U4162 ( .IN(n4516), .Q(n4665) );
  NBUFFX2 U4163 ( .IN(n4518), .Q(n4668) );
  NBUFFX2 U4164 ( .IN(n4363), .Q(n4674) );
  NBUFFX2 U4165 ( .IN(n4499), .Q(n4677) );
  NBUFFX2 U4166 ( .IN(n4520), .Q(n4678) );
  NBUFFX2 U4167 ( .IN(n4509), .Q(n4663) );
  NBUFFX2 U4168 ( .IN(n4511), .Q(n4666) );
  NBUFFX2 U4169 ( .IN(n4381), .Q(n4670) );
  NBUFFX2 U4170 ( .IN(n4506), .Q(n4675) );
  AOI21X1 U4171 ( .IN1(n2966), .IN2(n2672), .IN3(n2777), .QN(n2964) );
  NAND3X0 U4172 ( .IN1(n2968), .IN2(n2100), .IN3(n2829), .QN(n2966) );
  AOI21X1 U4173 ( .IN1(n2970), .IN2(n2687), .IN3(n2596), .QN(n2965) );
  NAND3X0 U4174 ( .IN1(n2972), .IN2(n1998), .IN3(n2839), .QN(n2970) );
  AOI21X1 U4175 ( .IN1(n2974), .IN2(n2754), .IN3(n2617), .QN(n2969) );
  NAND3X0 U4176 ( .IN1(n2976), .IN2(n1896), .IN3(n2809), .QN(n2974) );
  AOI21X1 U4177 ( .IN1(n2977), .IN2(n4498), .IN3(n2637), .QN(n2973) );
  NAND3X0 U4178 ( .IN1(n2979), .IN2(n1792), .IN3(n2819), .QN(n2977) );
  NAND2X0 U4179 ( .IN1(n2150), .IN2(n4660), .QN(n2351) );
  NAND2X0 U4180 ( .IN1(n2048), .IN2(n4658), .QN(n2279) );
  NAND2X0 U4181 ( .IN1(n1946), .IN2(n4656), .QN(n2207) );
  NAND2X0 U4182 ( .IN1(n1845), .IN2(n4654), .QN(n2430) );
  OA21X1 U4183 ( .IN1(n2793), .IN2(n1695), .IN3(n2095), .Q(n2780) );
  INVX0 U4184 ( .IN(n2794), .QN(n1695) );
  NOR3X0 U4185 ( .IN1(n2795), .IN2(n1690), .IN3(n2098), .QN(n2793) );
  INVX0 U4186 ( .IN(n2789), .QN(n1690) );
  OA21X1 U4187 ( .IN1(n2612), .IN2(n1638), .IN3(n1993), .Q(n2599) );
  INVX0 U4188 ( .IN(n2613), .QN(n1638) );
  NOR3X0 U4189 ( .IN1(n2614), .IN2(n1633), .IN3(n1996), .QN(n2612) );
  INVX0 U4190 ( .IN(n2608), .QN(n1633) );
  OA21X1 U4191 ( .IN1(n2633), .IN2(n1657), .IN3(n1891), .Q(n2620) );
  INVX0 U4192 ( .IN(n2634), .QN(n1657) );
  NOR3X0 U4193 ( .IN1(n2635), .IN2(n1652), .IN3(n1894), .QN(n2633) );
  INVX0 U4194 ( .IN(n2629), .QN(n1652) );
  NAND2X0 U4195 ( .IN1(n2150), .IN2(n4659), .QN(n2381) );
  NAND2X0 U4196 ( .IN1(n2048), .IN2(n4657), .QN(n2309) );
  NAND2X0 U4197 ( .IN1(n1946), .IN2(n4655), .QN(n2237) );
  NAND2X0 U4198 ( .IN1(n1845), .IN2(n4653), .QN(n2459) );
  NAND2X0 U4199 ( .IN1(n2790), .IN2(n2107), .QN(n2788) );
  NAND2X0 U4200 ( .IN1(n2609), .IN2(n2005), .QN(n2607) );
  NAND2X0 U4201 ( .IN1(n2630), .IN2(n1903), .QN(n2628) );
  NAND2X0 U4202 ( .IN1(n2650), .IN2(n1799), .QN(n2648) );
  NAND2X0 U4203 ( .IN1(n2795), .IN2(n2098), .QN(n2826) );
  NAND2X0 U4204 ( .IN1(n2614), .IN2(n1996), .QN(n2836) );
  NAND2X0 U4205 ( .IN1(n2635), .IN2(n1894), .QN(n2806) );
  NAND2X0 U4206 ( .IN1(n2655), .IN2(n1790), .QN(n2816) );
  INVX0 U4207 ( .IN(n2451), .QN(n1845) );
  INVX0 U4208 ( .IN(n2388), .QN(n2150) );
  INVX0 U4209 ( .IN(n2316), .QN(n2048) );
  INVX0 U4210 ( .IN(n2244), .QN(n1946) );
  INVX0 U4211 ( .IN(n2803), .QN(n1895) );
  OAI21X1 U4212 ( .IN1(n3269), .IN2(n2119), .IN3(n3267), .QN(n3278) );
  INVX0 U4213 ( .IN(n2968), .QN(n2096) );
  INVX0 U4214 ( .IN(n2972), .QN(n1994) );
  INVX0 U4215 ( .IN(n2976), .QN(n1892) );
  INVX0 U4216 ( .IN(n2979), .QN(n1788) );
  NAND2X0 U4217 ( .IN1(n1687), .IN2(n2107), .QN(n2792) );
  NAND2X0 U4218 ( .IN1(n1630), .IN2(n2005), .QN(n2611) );
  NAND2X0 U4219 ( .IN1(n1649), .IN2(n1903), .QN(n2632) );
  NAND2X0 U4220 ( .IN1(n1668), .IN2(n1799), .QN(n2652) );
  OA21X1 U4221 ( .IN1(n2653), .IN2(n1676), .IN3(n1787), .Q(n2640) );
  INVX0 U4222 ( .IN(n2654), .QN(n1676) );
  NOR3X0 U4223 ( .IN1(n2655), .IN2(n1671), .IN3(n1790), .QN(n2653) );
  INVX0 U4224 ( .IN(n2649), .QN(n1671) );
  NAND2X0 U4225 ( .IN1(n1607), .IN2(n2088), .QN(n3157) );
  NAND2X0 U4226 ( .IN1(n1986), .IN2(n1607), .QN(n3161) );
  NAND2X0 U4227 ( .IN1(n1884), .IN2(n1607), .QN(n3165) );
  NAND2X0 U4228 ( .IN1(n1780), .IN2(n1607), .QN(n3169) );
  NAND2X0 U4229 ( .IN1(n3196), .IN2(n3195), .QN(n3185) );
  NAND2X0 U4230 ( .IN1(n3212), .IN2(n3211), .QN(n3201) );
  NAND2X0 U4231 ( .IN1(n3225), .IN2(n3224), .QN(n3217) );
  NAND2X0 U4232 ( .IN1(n3237), .IN2(n3236), .QN(n3231) );
  OA21X1 U4233 ( .IN1(n4651), .IN2(n2097), .IN3(n2504), .Q(n3569) );
  OA21X1 U4234 ( .IN1(n4651), .IN2(n1995), .IN3(n2531), .Q(n3605) );
  OA21X1 U4235 ( .IN1(n4651), .IN2(n1893), .IN3(n2557), .Q(n3639) );
  OA21X1 U4236 ( .IN1(n4651), .IN2(n1789), .IN3(n2583), .Q(n3666) );
  INVX0 U4237 ( .IN(n4699), .QN(n4732) );
  AND4X1 U4238 ( .IN1(n3559), .IN2(n3535), .IN3(n3560), .IN4(n3520), .Q(n3522)
         );
  NAND2X0 U4239 ( .IN1(n4743), .IN2(n2127), .QN(n3559) );
  OA22X1_S38584 U4240 ( .IN1(n2127), .IN2(n3561), .IN3(n4743), .IN4(n3537), .Q(n3560)
         );
  INVX0 U4241 ( .IN(n4767), .QN(n4743) );
  AND4X1 U4242 ( .IN1(n3595), .IN2(n3570), .IN3(n3596), .IN4(n3546), .Q(n3548)
         );
  NAND2X0 U4243 ( .IN1(n4744), .IN2(n2025), .QN(n3595) );
  OA22X1_S38584 U4244 ( .IN1(n2025), .IN2(n3597), .IN3(n4745), .IN4(n3572), .Q(n3596)
         );
  NAND2X0 U4245 ( .IN1(n2029), .IN2(n4734), .QN(n3597) );
  AND4X1 U4246 ( .IN1(n3629), .IN2(n3606), .IN3(n3630), .IN4(n3581), .Q(n3583)
         );
  NAND2X0 U4247 ( .IN1(n4739), .IN2(n1923), .QN(n3629) );
  OA22X1_S38584 U4248 ( .IN1(n1923), .IN2(n3631), .IN3(n4747), .IN4(n3608), .Q(n3630)
         );
  NAND2X0 U4249 ( .IN1(n1927), .IN2(n4735), .QN(n3631) );
  AND4X1 U4250 ( .IN1(n3656), .IN2(n3640), .IN3(n3657), .IN4(n3617), .Q(n3619)
         );
  NAND2X0 U4251 ( .IN1(n4739), .IN2(n1821), .QN(n3656) );
  OA22X1_S38584 U4252 ( .IN1(n1821), .IN2(n3658), .IN3(n4750), .IN4(n3642), .Q(n3657)
         );
  NAND2X0 U4253 ( .IN1(n1825), .IN2(n4735), .QN(n3658) );
  INVX0 U4254 ( .IN(n4699), .QN(n4733) );
  INVX0 U4255 ( .IN(g26135), .QN(n1575) );
  INVX0 U4256 ( .IN(n4770), .QN(n4738) );
  INVX0 U4257 ( .IN(n4771), .QN(n4770) );
  INVX0 U4258 ( .IN(n4772), .QN(n4767) );
  INVX0 U4259 ( .IN(n4772), .QN(n4768) );
  INVX0 U4260 ( .IN(n4773), .QN(n4765) );
  INVX0 U4261 ( .IN(n4772), .QN(n4766) );
  INVX0 U4262 ( .IN(n4773), .QN(n4764) );
  INVX0 U4263 ( .IN(n4775), .QN(n4760) );
  INVX0 U4264 ( .IN(n4771), .QN(n4769) );
  INVX0 U4265 ( .IN(n4775), .QN(n4761) );
  INVX0 U4266 ( .IN(n4728), .QN(n4721) );
  INVX0 U4267 ( .IN(n4728), .QN(n4720) );
  INVX0 U4268 ( .IN(n4716), .QN(n4717) );
  INVX0 U4269 ( .IN(n4729), .QN(n4718) );
  INVX0 U4270 ( .IN(n4729), .QN(n4719) );
  INVX0 U4271 ( .IN(n4727), .QN(n4722) );
  INVX0 U4272 ( .IN(n4727), .QN(n4723) );
  INVX0 U4273 ( .IN(n4724), .QN(n4700) );
  INVX0 U4274 ( .IN(n4724), .QN(n4701) );
  NAND2X0 U4275 ( .IN1(n3186), .IN2(n3185), .QN(n3178) );
  NAND2X0 U4276 ( .IN1(n3202), .IN2(n3201), .QN(n3183) );
  NAND2X0 U4277 ( .IN1(n3218), .IN2(n3217), .QN(n3191) );
  NAND2X0 U4278 ( .IN1(n3232), .IN2(n3231), .QN(n3207) );
  NOR2X0 U4279 ( .IN1(n2131), .IN2(n4734), .QN(n3509) );
  NOR2X0 U4280 ( .IN1(n2104), .IN2(n4734), .QN(n3539) );
  NOR2X0 U4281 ( .IN1(n2029), .IN2(n4734), .QN(n3526) );
  NOR2X0 U4282 ( .IN1(n2002), .IN2(n4734), .QN(n3574) );
  NOR2X0 U4283 ( .IN1(n1927), .IN2(n4734), .QN(n3552) );
  NOR2X0 U4284 ( .IN1(n1900), .IN2(n4734), .QN(n3610) );
  NOR2X0 U4285 ( .IN1(n1825), .IN2(n4734), .QN(n3587) );
  NOR2X0 U4286 ( .IN1(n1796), .IN2(n4734), .QN(n3644) );
  AO21X1 U4287 ( .IN1(n2017), .IN2(n3322), .IN3(n2015), .Q(n3321) );
  NAND2X0 U4288 ( .IN1(n2016), .IN2(n2027), .QN(n3322) );
  INVX0 U4289 ( .IN(n3323), .QN(n2015) );
  AO21X1 U4290 ( .IN1(n1915), .IN2(n3362), .IN3(n1913), .Q(n3361) );
  NAND2X0 U4291 ( .IN1(n1914), .IN2(n1925), .QN(n3362) );
  INVX0 U4292 ( .IN(n3363), .QN(n1913) );
  AO21X1 U4293 ( .IN1(n1811), .IN2(n3401), .IN3(n1809), .Q(n3400) );
  NAND2X0 U4294 ( .IN1(n1810), .IN2(n1823), .QN(n3401) );
  INVX0 U4295 ( .IN(n3402), .QN(n1809) );
  NAND3X0 U4296 ( .IN1(n4759), .IN2(n2131), .IN3(n2128), .QN(n3520) );
  NAND3X0 U4297 ( .IN1(n4759), .IN2(n2029), .IN3(n2026), .QN(n3546) );
  NAND3X0 U4298 ( .IN1(n4758), .IN2(n1927), .IN3(n1924), .QN(n3581) );
  NAND3X0 U4299 ( .IN1(n4758), .IN2(n1825), .IN3(n1822), .QN(n3617) );
  NAND3X0 U4300 ( .IN1(n2129), .IN2(n2131), .IN3(n4757), .QN(n3535) );
  NAND3X0 U4301 ( .IN1(n2027), .IN2(n2029), .IN3(n4755), .QN(n3570) );
  NAND3X0 U4302 ( .IN1(n1925), .IN2(n1927), .IN3(n4754), .QN(n3606) );
  NAND3X0 U4303 ( .IN1(n1823), .IN2(n1825), .IN3(n4756), .QN(n3640) );
  NAND3X0 U4304 ( .IN1(n2103), .IN2(n2104), .IN3(n4755), .QN(n3592) );
  NAND3X0 U4305 ( .IN1(n2001), .IN2(n2002), .IN3(n4755), .QN(n3626) );
  NAND3X0 U4306 ( .IN1(n1899), .IN2(n1900), .IN3(n4756), .QN(n3653) );
  NAND3X0 U4307 ( .IN1(n1795), .IN2(n1796), .IN3(n4756), .QN(n3671) );
  NAND2X0 U4308 ( .IN1(n3936), .IN2(n1748), .QN(n3906) );
  NAND2X0 U4309 ( .IN1(n2131), .IN2(n4734), .QN(n3561) );
  NAND2X0 U4310 ( .IN1(n2104), .IN2(n4735), .QN(n3624) );
  NAND2X0 U4311 ( .IN1(n2002), .IN2(n4735), .QN(n3651) );
  NAND2X0 U4312 ( .IN1(n1900), .IN2(n4735), .QN(n3669) );
  NAND2X0 U4313 ( .IN1(n1796), .IN2(n4735), .QN(n3676) );
  INVX0 U4314 ( .IN(n3734), .QN(n1586) );
  INVX0 U4315 ( .IN(n4031), .QN(n1590) );
  INVX0 U4316 ( .IN(n4032), .QN(n1591) );
  INVX0 U4317 ( .IN(n4034), .QN(n1593) );
  INVX0 U4318 ( .IN(n4033), .QN(n1592) );
  INVX0 U4319 ( .IN(n4037), .QN(n1594) );
  INVX0 U4320 ( .IN(n4040), .QN(n1596) );
  INVX0 U4321 ( .IN(n4038), .QN(n1595) );
  INVX0 U4322 ( .IN(n4043), .QN(n1597) );
  INVX0 U4323 ( .IN(n4046), .QN(n1599) );
  INVX0 U4324 ( .IN(n4044), .QN(n1598) );
  INVX0 U4325 ( .IN(n4049), .QN(n1600) );
  INVX0 U4326 ( .IN(n4051), .QN(n1601) );
  INVX0 U4327 ( .IN(n2490), .QN(n2097) );
  INVX0 U4328 ( .IN(n2517), .QN(n1995) );
  INVX0 U4329 ( .IN(n2543), .QN(n1893) );
  INVX0 U4330 ( .IN(n2569), .QN(n1789) );
  OAI21X1 U4331 ( .IN1(n3310), .IN2(n2017), .IN3(n3308), .QN(n3319) );
  OAI21X1 U4332 ( .IN1(n3350), .IN2(n1915), .IN3(n3348), .QN(n3359) );
  OAI21X1 U4333 ( .IN1(n3389), .IN2(n1811), .IN3(n3387), .QN(n3398) );
  INVX0 U4334 ( .IN(n3698), .QN(n1745) );
  INVX0 U4335 ( .IN(n3513), .QN(n1619) );
  INVX0 U4336 ( .IN(n3523), .QN(n1618) );
  INVX0 U4337 ( .IN(n3538), .QN(n1617) );
  INVX0 U4338 ( .IN(n3530), .QN(n1616) );
  INVX0 U4339 ( .IN(n3549), .QN(n1615) );
  INVX0 U4340 ( .IN(n3573), .QN(n1614) );
  INVX0 U4341 ( .IN(n3556), .QN(n1613) );
  INVX0 U4342 ( .IN(n3584), .QN(n1612) );
  INVX0 U4343 ( .IN(n3609), .QN(n1611) );
  INVX0 U4344 ( .IN(n3591), .QN(n1610) );
  INVX0 U4345 ( .IN(n3620), .QN(n1609) );
  INVX0 U4346 ( .IN(n3643), .QN(n1608) );
  NAND2X0 U4347 ( .IN1(n2106), .IN2(n1693), .QN(n3002) );
  NAND2X0 U4348 ( .IN1(n2004), .IN2(n1636), .QN(n3010) );
  NAND2X0 U4349 ( .IN1(n1798), .IN2(n1674), .QN(n3025) );
  NAND2X0 U4350 ( .IN1(n1902), .IN2(n1655), .QN(n3018) );
  INVX0 U4351 ( .IN(n3186), .QN(n2089) );
  INVX0 U4352 ( .IN(n3202), .QN(n1987) );
  INVX0 U4353 ( .IN(n3218), .QN(n1885) );
  INVX0 U4354 ( .IN(n3232), .QN(n1781) );
  INVX0 U4355 ( .IN(n3916), .QN(n1746) );
  INVX0 U4356 ( .IN(n3290), .QN(n2128) );
  INVX0 U4357 ( .IN(n3331), .QN(n2026) );
  INVX0 U4358 ( .IN(n3371), .QN(n1924) );
  INVX0 U4359 ( .IN(n3410), .QN(n1822) );
  INVX0 U4360 ( .IN(n3197), .QN(n1693) );
  INVX0 U4361 ( .IN(n3213), .QN(n1636) );
  INVX0 U4362 ( .IN(n3226), .QN(n1655) );
  INVX0 U4363 ( .IN(n3238), .QN(n1674) );
  INVX0 U4364 ( .IN(n4651), .QN(n1607) );
  INVX0 U4365 ( .IN(n2504), .QN(n2092) );
  INVX0 U4366 ( .IN(n2531), .QN(n1990) );
  INVX0 U4367 ( .IN(n2557), .QN(n1888) );
  INVX0 U4368 ( .IN(n2583), .QN(n1784) );
  AO221X1 U4369 ( .IN1(n2456), .IN2(n4653), .IN3(n2438), .IN4(n1852), .IN5(
        n2439), .Q(n2417) );
  AOI221X1 U4370 ( .IN1(n2442), .IN2(n4654), .IN3(n2433), .IN4(n1847), .IN5(
        n2439), .QN(n2413) );
  AOI221X1 U4371 ( .IN1(n2448), .IN2(n4654), .IN3(n2433), .IN4(n1850), .IN5(
        n2439), .QN(n2418) );
  AOI221X1 U4372 ( .IN1(n2444), .IN2(n4653), .IN3(n2438), .IN4(n1849), .IN5(
        n2439), .QN(n2412) );
  NOR2X0 U4373 ( .IN1(n2365), .IN2(n2136), .QN(n2361) );
  NOR2X0 U4374 ( .IN1(n2221), .IN2(n1932), .QN(n2217) );
  NAND2X0 U4375 ( .IN1(n2478), .IN2(n2453), .QN(n2454) );
  AND4X1 U4376 ( .IN1(n1584), .IN2(n2469), .IN3(n2470), .IN4(n2459), .Q(n2414)
         );
  NAND2X0 U4377 ( .IN1(n2471), .IN2(n4653), .QN(n2470) );
  NAND2X0 U4378 ( .IN1(n2438), .IN2(n1855), .QN(n2469) );
  AND4X1 U4379 ( .IN1(n1584), .IN2(n2428), .IN3(n2429), .IN4(n2430), .Q(n2411)
         );
  NAND2X0 U4380 ( .IN1(n2431), .IN2(n4654), .QN(n2429) );
  NAND2X0 U4381 ( .IN1(n2433), .IN2(n1851), .QN(n2428) );
  NAND4X0 U4382 ( .IN1(n1584), .IN2(n2457), .IN3(n2458), .IN4(n2459), .QN(
        n2405) );
  NAND2X0 U4383 ( .IN1(n2460), .IN2(n4653), .QN(n2458) );
  NAND2X0 U4384 ( .IN1(n2438), .IN2(n1846), .QN(n2457) );
  NAND4X0 U4385 ( .IN1(n1584), .IN2(n2462), .IN3(n2463), .IN4(n2430), .QN(
        n2416) );
  NAND2X0 U4386 ( .IN1(n2464), .IN2(n4654), .QN(n2463) );
  NAND2X0 U4387 ( .IN1(n2433), .IN2(n1854), .QN(n2462) );
  NAND4X0 U4388 ( .IN1(n1584), .IN2(n2465), .IN3(n2466), .IN4(n2430), .QN(
        n2404) );
  NAND2X0 U4389 ( .IN1(n2467), .IN2(n4654), .QN(n2466) );
  NAND2X0 U4390 ( .IN1(n2433), .IN2(n1848), .QN(n2465) );
  AOI221X1 U4391 ( .IN1(n2436), .IN2(n4653), .IN3(n2438), .IN4(n1853), .IN5(
        n2439), .QN(n2409) );
  INVX0 U4392 ( .IN(n2453), .QN(n1832) );
  XOR2X1 U4393 ( .IN1(n2502), .IN2(n2672), .Q(n2735) );
  XOR2X1 U4394 ( .IN1(n2529), .IN2(n2687), .Q(n2750) );
  XOR2X1 U4395 ( .IN1(n2581), .IN2(n4498), .Q(n2774) );
  NAND2X0 U4396 ( .IN1(n2361), .IN2(n2374), .QN(n2355) );
  NAND2X0 U4397 ( .IN1(n2289), .IN2(n2302), .QN(n2283) );
  NAND2X0 U4398 ( .IN1(n2217), .IN2(n2230), .QN(n2211) );
  NAND2X0 U4399 ( .IN1(n2446), .IN2(n2445), .QN(n2434) );
  NAND2X0 U4400 ( .IN1(n2385), .IN2(n2363), .QN(n2364) );
  NAND2X0 U4401 ( .IN1(n2424), .IN2(n1582), .QN(n3740) );
  AO22X1 U4402 ( .IN1(n4136), .IN2(n2180), .IN3(n4137), .IN4(n2124), .Q(g22687) );
  INVX0 U4403 ( .IN(n3843), .QN(n2124) );
  NAND2X0 U4404 ( .IN1(n4660), .IN2(n3843), .QN(n4136) );
  NOR2X0 U4405 ( .IN1(n2126), .IN2(n4303), .QN(n4137) );
  AO22X1 U4406 ( .IN1(n4138), .IN2(n2180), .IN3(n4139), .IN4(n2022), .Q(g22651) );
  INVX0 U4407 ( .IN(n3845), .QN(n2022) );
  NAND2X0 U4408 ( .IN1(n4658), .IN2(n3845), .QN(n4138) );
  NOR2X0 U4409 ( .IN1(n2024), .IN2(n4297), .QN(n4139) );
  AO22X1 U4410 ( .IN1(n4140), .IN2(n2180), .IN3(n4141), .IN4(n1920), .Q(g22615) );
  INVX0 U4411 ( .IN(n3847), .QN(n1920) );
  NAND2X0 U4412 ( .IN1(n4656), .IN2(n3847), .QN(n4140) );
  NOR2X0 U4413 ( .IN1(n1922), .IN2(n4304), .QN(n4141) );
  AO22X1 U4414 ( .IN1(n4142), .IN2(n2180), .IN3(n4143), .IN4(n1816), .Q(g22578) );
  INVX0 U4415 ( .IN(n3848), .QN(n1816) );
  NAND2X0 U4416 ( .IN1(n4654), .IN2(n3848), .QN(n4142) );
  NOR2X0 U4417 ( .IN1(n1820), .IN2(n4310), .QN(n4143) );
  NAND2X0 U4418 ( .IN1(n2778), .IN2(n2099), .QN(n2490) );
  NAND2X0 U4419 ( .IN1(n2597), .IN2(n1997), .QN(n2517) );
  NAND2X0 U4420 ( .IN1(n2638), .IN2(n1791), .QN(n2569) );
  NAND2X0 U4421 ( .IN1(n4599), .IN2(g22687), .QN(n3503) );
  NAND2X0 U4422 ( .IN1(n4602), .IN2(g22687), .QN(n3504) );
  NAND2X0 U4423 ( .IN1(g7302), .IN2(g22687), .QN(n3508) );
  NAND2X0 U4424 ( .IN1(n4611), .IN2(g22651), .QN(n3507) );
  NAND2X0 U4425 ( .IN1(n4614), .IN2(g22651), .QN(n3514) );
  NAND2X0 U4426 ( .IN1(g7052), .IN2(g22651), .QN(n3525) );
  NAND2X0 U4427 ( .IN1(n4623), .IN2(g22615), .QN(n3517) );
  NAND2X0 U4428 ( .IN1(n4626), .IN2(g22615), .QN(n3531) );
  NAND2X0 U4429 ( .IN1(g6750), .IN2(g22615), .QN(n3551) );
  NAND2X0 U4430 ( .IN1(n4633), .IN2(g22578), .QN(n3534) );
  NAND2X0 U4431 ( .IN1(n4636), .IN2(g22578), .QN(n3557) );
  NAND2X0 U4432 ( .IN1(g6485), .IN2(g22578), .QN(n3586) );
  AND3X1 U4433 ( .IN1(n2710), .IN2(n2905), .IN3(n2663), .Q(n2843) );
  XOR2X1 U4434 ( .IN1(n2708), .IN2(n2672), .Q(n2905) );
  AND3X1 U4435 ( .IN1(n2729), .IN2(n2923), .IN3(n2677), .Q(n2848) );
  XOR2X1 U4436 ( .IN1(n2727), .IN2(n2687), .Q(n2923) );
  AND3X1 U4437 ( .IN1(n2761), .IN2(n2958), .IN3(n2706), .Q(n2863) );
  XOR2X1 U4438 ( .IN1(n2759), .IN2(n4498), .Q(n2958) );
  AND3X1 U4439 ( .IN1(n2867), .IN2(n2904), .IN3(n2843), .Q(n2736) );
  XOR2X1 U4440 ( .IN1(n2503), .IN2(n2672), .Q(n2904) );
  AND3X1 U4441 ( .IN1(n2875), .IN2(n2922), .IN3(n2848), .Q(n2751) );
  XOR2X1 U4442 ( .IN1(n2530), .IN2(n2687), .Q(n2922) );
  AND3X1 U4443 ( .IN1(n2889), .IN2(n2957), .IN3(n2863), .Q(n2775) );
  XOR2X1 U4444 ( .IN1(n2582), .IN2(n4498), .Q(n2957) );
  AND3X1 U4445 ( .IN1(n2906), .IN2(n2725), .IN3(n2724), .Q(n2663) );
  XOR2X1 U4446 ( .IN1(n2512), .IN2(n2672), .Q(n2906) );
  AND3X1 U4447 ( .IN1(n2924), .IN2(n2741), .IN3(n2740), .Q(n2677) );
  XOR2X1 U4448 ( .IN1(n2538), .IN2(n2687), .Q(n2924) );
  AND3X1 U4449 ( .IN1(n2959), .IN2(n2771), .IN3(n2770), .Q(n2706) );
  XOR2X1 U4450 ( .IN1(n2590), .IN2(n2720), .Q(n2959) );
  NOR4X0 U4451 ( .IN1(n2476), .IN2(n1847), .IN3(n1850), .IN4(n1849), .QN(n2472) );
  NOR4X0 U4452 ( .IN1(n2474), .IN2(n2467), .IN3(n2475), .IN4(n2460), .QN(n2473) );
  NAND3X0 U4453 ( .IN1(n2456), .IN2(n2477), .IN3(n2436), .QN(n2476) );
  NOR4X0 U4454 ( .IN1(n2398), .IN2(n2152), .IN3(n2155), .IN4(n2154), .QN(n2394) );
  NOR4X0 U4455 ( .IN1(n2396), .IN2(n2371), .IN3(n2397), .IN4(n2393), .QN(n2395) );
  NAND3X0 U4456 ( .IN1(n2390), .IN2(n2399), .IN3(n2357), .QN(n2398) );
  NOR4X0 U4457 ( .IN1(n2326), .IN2(n2050), .IN3(n2053), .IN4(n2052), .QN(n2322) );
  NOR4X0 U4458 ( .IN1(n2324), .IN2(n2299), .IN3(n2325), .IN4(n2321), .QN(n2323) );
  NAND3X0 U4459 ( .IN1(n2318), .IN2(n2327), .IN3(n2285), .QN(n2326) );
  NOR4X0 U4460 ( .IN1(n2254), .IN2(n1948), .IN3(n1951), .IN4(n1950), .QN(n2250) );
  NOR4X0 U4461 ( .IN1(n2252), .IN2(n2227), .IN3(n2253), .IN4(n2249), .QN(n2251) );
  NAND3X0 U4462 ( .IN1(n2246), .IN2(n2255), .IN3(n2213), .QN(n2254) );
  AO22X1 U4463 ( .IN1(n4662), .IN2(n4660), .IN3(n3260), .IN4(n3255), .Q(n3249)
         );
  NOR2X0 U4464 ( .IN1(n3283), .IN2(n4662), .QN(n3260) );
  OA22X1_S38584 U4465 ( .IN1(n1765), .IN2(n3256), .IN3(n3253), .IN4(n3257), .Q(n3283)
         );
  AO22X1 U4466 ( .IN1(n4661), .IN2(n4659), .IN3(n3252), .IN4(n4553), .Q(n3248)
         );
  ISOLANDX1 U4467 ( .D(n3253), .ISO(n3254), .Q(n3252) );
  OA22X1_S38584 U4468 ( .IN1(n3255), .IN2(n3256), .IN3(n1766), .IN4(n3257), .Q(n3254)
         );
  AO22X1 U4469 ( .IN1(n4661), .IN2(n4658), .IN3(n3301), .IN4(n3296), .Q(n3258)
         );
  NOR2X0 U4470 ( .IN1(n3324), .IN2(n4661), .QN(n3301) );
  OA22X1_S38584 U4471 ( .IN1(n1763), .IN2(n3297), .IN3(n3294), .IN4(n3298), .Q(n3324)
         );
  AO22X1 U4472 ( .IN1(n4662), .IN2(n4657), .IN3(n3293), .IN4(n3294), .Q(n3250)
         );
  NOR2X0 U4473 ( .IN1(n3295), .IN2(n4662), .QN(n3293) );
  OA22X1_S38584 U4474 ( .IN1(n3296), .IN2(n3297), .IN3(n1764), .IN4(n3298), .Q(n3295)
         );
  AO22X1 U4475 ( .IN1(n4661), .IN2(n4656), .IN3(n3341), .IN4(n3337), .Q(n3299)
         );
  NOR2X0 U4476 ( .IN1(n3364), .IN2(n4661), .QN(n3341) );
  OA22X1_S38584 U4477 ( .IN1(n1761), .IN2(n3338), .IN3(n3335), .IN4(n3339), .Q(n3364)
         );
  AO22X1 U4478 ( .IN1(n4661), .IN2(n4655), .IN3(n3334), .IN4(n3335), .Q(n3259)
         );
  NOR2X0 U4479 ( .IN1(n3336), .IN2(n4661), .QN(n3334) );
  OA22X1_S38584 U4480 ( .IN1(n3337), .IN2(n3338), .IN3(n1762), .IN4(n3339), .Q(n3336)
         );
  AO22X1 U4481 ( .IN1(n4662), .IN2(n4654), .IN3(n3380), .IN4(n3377), .Q(n3340)
         );
  NOR2X0 U4482 ( .IN1(n3403), .IN2(n4661), .QN(n3380) );
  OA22X1_S38584 U4483 ( .IN1(n1759), .IN2(n3378), .IN3(n3375), .IN4(n3379), .Q(n3403)
         );
  AND4X1 U4484 ( .IN1(n1569), .IN2(n2379), .IN3(n2380), .IN4(n2381), .Q(n2342)
         );
  NAND2X0 U4485 ( .IN1(n2382), .IN2(n4659), .QN(n2380) );
  NAND2X0 U4486 ( .IN1(n2359), .IN2(n2160), .QN(n2379) );
  AND4X1 U4487 ( .IN1(n1567), .IN2(n2307), .IN3(n2308), .IN4(n2309), .Q(n2270)
         );
  NAND2X0 U4488 ( .IN1(n2310), .IN2(n4657), .QN(n2308) );
  NAND2X0 U4489 ( .IN1(n2287), .IN2(n2058), .QN(n2307) );
  AND4X1 U4490 ( .IN1(n1569), .IN2(n2349), .IN3(n2350), .IN4(n2351), .Q(n2339)
         );
  NAND2X0 U4491 ( .IN1(n2352), .IN2(n4660), .QN(n2350) );
  NAND2X0 U4492 ( .IN1(n2354), .IN2(n2156), .QN(n2349) );
  AND4X1 U4493 ( .IN1(n1567), .IN2(n2277), .IN3(n2278), .IN4(n2279), .Q(n2267)
         );
  NAND2X0 U4494 ( .IN1(n2280), .IN2(n4658), .QN(n2278) );
  NAND2X0 U4495 ( .IN1(n2282), .IN2(n2054), .QN(n2277) );
  AO221X1 U4496 ( .IN1(n2390), .IN2(n4659), .IN3(n2359), .IN4(n2157), .IN5(
        n2360), .Q(n2345) );
  AO221X1 U4497 ( .IN1(n2318), .IN2(n4657), .IN3(n2287), .IN4(n2055), .IN5(
        n2288), .Q(n2273) );
  AO221X1 U4498 ( .IN1(n2246), .IN2(n4655), .IN3(n2215), .IN4(n1953), .IN5(
        n2216), .Q(n2201) );
  INVX0 U4499 ( .IN(n2288), .QN(n1567) );
  NOR2X0 U4500 ( .IN1(n4481), .IN2(n2424), .QN(n2425) );
  NAND2X0 U4501 ( .IN1(n4597), .IN2(n4129), .QN(n2424) );
  XOR2X1 U4502 ( .IN1(n2672), .IN2(n2501), .Q(n2734) );
  XOR2X1 U4503 ( .IN1(n2687), .IN2(n2528), .Q(n2749) );
  XOR2X1 U4504 ( .IN1(n4498), .IN2(n2580), .Q(n2773) );
  XOR2X1 U4505 ( .IN1(n4508), .IN2(n2511), .Q(n2867) );
  XOR2X1 U4506 ( .IN1(n4510), .IN2(n2537), .Q(n2875) );
  XOR2X1 U4507 ( .IN1(n1785), .IN2(n2589), .Q(n2889) );
  NAND4X0 U4508 ( .IN1(n1569), .IN2(n2366), .IN3(n2367), .IN4(n2351), .QN(
        n2341) );
  NAND2X0 U4509 ( .IN1(n2368), .IN2(n4660), .QN(n2367) );
  NAND2X0 U4510 ( .IN1(n2354), .IN2(n2159), .QN(n2366) );
  NAND4X0 U4511 ( .IN1(n1567), .IN2(n2294), .IN3(n2295), .IN4(n2279), .QN(
        n2269) );
  NAND2X0 U4512 ( .IN1(n2296), .IN2(n4658), .QN(n2295) );
  NAND2X0 U4513 ( .IN1(n2282), .IN2(n2057), .QN(n2294) );
  NAND4X0 U4514 ( .IN1(n1565), .IN2(n2222), .IN3(n2223), .IN4(n2207), .QN(
        n2197) );
  NAND2X0 U4515 ( .IN1(n2224), .IN2(n4656), .QN(n2223) );
  NAND2X0 U4516 ( .IN1(n2210), .IN2(n1955), .QN(n2222) );
  NAND4X0 U4517 ( .IN1(n1569), .IN2(n2369), .IN3(n2370), .IN4(n2351), .QN(
        n2333) );
  NAND2X0 U4518 ( .IN1(n2371), .IN2(n4660), .QN(n2370) );
  NAND2X0 U4519 ( .IN1(n2354), .IN2(n2153), .QN(n2369) );
  NAND4X0 U4520 ( .IN1(n1569), .IN2(n2391), .IN3(n2392), .IN4(n2381), .QN(
        n2332) );
  NAND2X0 U4521 ( .IN1(n2393), .IN2(n4659), .QN(n2392) );
  NAND2X0 U4522 ( .IN1(n2359), .IN2(n2151), .QN(n2391) );
  NAND2X0 U4523 ( .IN1(n3740), .IN2(n1582), .QN(n3858) );
  NOR2X0 U4524 ( .IN1(n4480), .IN2(n4102), .QN(n4056) );
  AOI221X1 U4525 ( .IN1(n2659), .IN2(n2666), .IN3(n2661), .IN4(n2667), .IN5(
        n2668), .QN(n2657) );
  XNOR2X1 U4526 ( .IN1(n2499), .IN2(n2669), .Q(n2667) );
  XOR2X1 U4527 ( .IN1(n2500), .IN2(n2672), .Q(n2671) );
  AOI221X1 U4528 ( .IN1(n2673), .IN2(n2681), .IN3(n2675), .IN4(n2682), .IN5(
        n2683), .QN(n2664) );
  XNOR2X1 U4529 ( .IN1(n2526), .IN2(n2684), .Q(n2682) );
  XOR2X1 U4530 ( .IN1(n2527), .IN2(n2687), .Q(n2686) );
  AOI221X1 U4531 ( .IN1(n2702), .IN2(n2714), .IN3(n2704), .IN4(n2715), .IN5(
        n2716), .QN(n2693) );
  XNOR2X1 U4532 ( .IN1(n2578), .IN2(n2717), .Q(n2715) );
  XOR2X1 U4533 ( .IN1(n2579), .IN2(n4498), .Q(n2719) );
  INVX0 U4534 ( .IN(n4144), .QN(n2180) );
  OA21X1 U4535 ( .IN1(n3740), .IN2(n3857), .IN3(n3858), .Q(g26048) );
  XOR2X1 U4536 ( .IN1(n4354), .IN2(n3859), .Q(n3857) );
  INVX0 U4537 ( .IN(n4362), .QN(n4689) );
  AOI221X1 U4538 ( .IN1(n2384), .IN2(n4659), .IN3(n2359), .IN4(n2154), .IN5(
        n2360), .QN(n2346) );
  AOI221X1 U4539 ( .IN1(n2312), .IN2(n4657), .IN3(n2287), .IN4(n2052), .IN5(
        n2288), .QN(n2274) );
  AOI221X1 U4540 ( .IN1(n2240), .IN2(n4655), .IN3(n2215), .IN4(n1950), .IN5(
        n2216), .QN(n2202) );
  AOI221X1 U4541 ( .IN1(n2357), .IN2(n4659), .IN3(n2359), .IN4(n2158), .IN5(
        n2360), .QN(n2337) );
  AOI221X1 U4542 ( .IN1(n2285), .IN2(n4657), .IN3(n2287), .IN4(n2056), .IN5(
        n2288), .QN(n2265) );
  AOI221X1 U4543 ( .IN1(n2373), .IN2(n4660), .IN3(n2354), .IN4(n2155), .IN5(
        n2360), .QN(n2340) );
  AOI221X1 U4544 ( .IN1(n2301), .IN2(n4658), .IN3(n2282), .IN4(n2053), .IN5(
        n2288), .QN(n2268) );
  AOI221X1 U4545 ( .IN1(n2229), .IN2(n4656), .IN3(n2210), .IN4(n1951), .IN5(
        n2216), .QN(n2196) );
  AOI221X1 U4546 ( .IN1(n2377), .IN2(n4660), .IN3(n2354), .IN4(n2152), .IN5(
        n2360), .QN(n2344) );
  AOI221X1 U4547 ( .IN1(n2305), .IN2(n4658), .IN3(n2282), .IN4(n2050), .IN5(
        n2288), .QN(n2272) );
  AO22X1 U4548 ( .IN1(n4662), .IN2(n4653), .IN3(n3374), .IN4(n3375), .Q(n3300)
         );
  NOR2X0 U4549 ( .IN1(n3376), .IN2(n4661), .QN(n3374) );
  OA22X1_S38584 U4550 ( .IN1(n3377), .IN2(n3378), .IN3(n1760), .IN4(n3379), .Q(n3376)
         );
  NAND2X0 U4551 ( .IN1(n2422), .IN2(n2423), .QN(n4262) );
  AO21X1 U4552 ( .IN1(n4481), .IN2(n2424), .IN3(n2425), .Q(n2423) );
  NOR2X0 U4553 ( .IN1(n1580), .IN2(n4120), .QN(g23359) );
  XOR2X1 U4554 ( .IN1(n2425), .IN2(n4350), .Q(n4120) );
  INVX0 U4555 ( .IN(n2422), .QN(n1580) );
  INVX0 U4556 ( .IN(n2961), .QN(n1818) );
  INVX0 U4557 ( .IN(n3156), .QN(n1817) );
  INVX0 U4558 ( .IN(n4553), .QN(n4662) );
  INVX0 U4559 ( .IN(n4553), .QN(n4661) );
  INVX0 U4560 ( .IN(n4514), .QN(n4587) );
  INVX0 U4561 ( .IN(n4515), .QN(n4589) );
  INVX0 U4562 ( .IN(n4512), .QN(n4593) );
  NAND2X0 U4563 ( .IN1(n2313), .IN2(n2291), .QN(n2292) );
  NAND2X0 U4564 ( .IN1(n2241), .IN2(n2219), .QN(n2220) );
  NAND4X0 U4565 ( .IN1(n3863), .IN2(n3864), .IN3(n3865), .IN4(n3866), .QN(
        n2899) );
  XNOR2X1 U4566 ( .IN1(n2666), .IN2(n3884), .Q(n3864) );
  XOR2X1 U4567 ( .IN1(n2081), .IN2(n3885), .Q(n3863) );
  NOR3X0 U4568 ( .IN1(n2082), .IN2(n3880), .IN3(n3881), .QN(n3865) );
  NAND4X0 U4569 ( .IN1(n3760), .IN2(n3761), .IN3(n3762), .IN4(n3763), .QN(
        n2917) );
  XNOR2X1 U4570 ( .IN1(n2681), .IN2(n3781), .Q(n3761) );
  XOR2X1 U4571 ( .IN1(n1979), .IN2(n3782), .Q(n3760) );
  NOR3X0 U4572 ( .IN1(n1980), .IN2(n3777), .IN3(n3778), .QN(n3762) );
  NAND4X0 U4573 ( .IN1(n3790), .IN2(n3791), .IN3(n3792), .IN4(n3793), .QN(
        n2935) );
  XNOR2X1 U4574 ( .IN1(n2696), .IN2(n3811), .Q(n3791) );
  XOR2X1 U4575 ( .IN1(n1877), .IN2(n3812), .Q(n3790) );
  NOR3X0 U4576 ( .IN1(n1878), .IN2(n3807), .IN3(n3808), .QN(n3792) );
  NAND4X0 U4577 ( .IN1(n3818), .IN2(n3819), .IN3(n3820), .IN4(n3821), .QN(
        n2952) );
  XNOR2X1 U4578 ( .IN1(n2714), .IN2(n3839), .Q(n3819) );
  XOR2X1 U4579 ( .IN1(n1773), .IN2(n3840), .Q(n3818) );
  NOR3X0 U4580 ( .IN1(n1774), .IN2(n3835), .IN3(n3836), .QN(n3820) );
  NAND2X0 U4581 ( .IN1(n2618), .IN2(n1895), .QN(n2543) );
  NAND2X0 U4582 ( .IN1(n2627), .IN2(n4118), .QN(n2803) );
  NOR2X0 U4583 ( .IN1(n2899), .IN2(n2967), .QN(n2777) );
  NOR2X0 U4584 ( .IN1(n2917), .IN2(n2971), .QN(n2596) );
  NOR2X0 U4585 ( .IN1(n2935), .IN2(n2975), .QN(n2617) );
  NOR2X0 U4586 ( .IN1(n2952), .IN2(n2978), .QN(n2637) );
  OA22X1_S38584 U4587 ( .IN1(n4385), .IN2(n2968), .IN3(n2795), .IN4(n2096), .Q(n3030)
         );
  OA22X1_S38584 U4588 ( .IN1(n4386), .IN2(n2972), .IN3(n2614), .IN4(n1994), .Q(n3034)
         );
  OA22X1_S38584 U4589 ( .IN1(n4387), .IN2(n2976), .IN3(n2635), .IN4(n1892), .Q(n3066)
         );
  OA22X1_S38584 U4590 ( .IN1(n4388), .IN2(n2979), .IN3(n2655), .IN4(n1788), .Q(n3098)
         );
  NAND2X0 U4591 ( .IN1(n3038), .IN2(n3050), .QN(n2789) );
  NAND3X0 U4592 ( .IN1(n3051), .IN2(n3052), .IN3(n3053), .QN(n3050) );
  AO221X1 U4593 ( .IN1(n3054), .IN2(n3057), .IN3(n3056), .IN4(n1697), .IN5(
        n3055), .Q(n3051) );
  NAND3X0 U4594 ( .IN1(n3058), .IN2(n3059), .IN3(n3060), .QN(n3052) );
  NAND2X0 U4595 ( .IN1(n3070), .IN2(n3082), .QN(n2608) );
  NAND3X0 U4596 ( .IN1(n3083), .IN2(n3084), .IN3(n3085), .QN(n3082) );
  AO221X1 U4597 ( .IN1(n3086), .IN2(n3089), .IN3(n3088), .IN4(n1640), .IN5(
        n3087), .Q(n3083) );
  NAND3X0 U4598 ( .IN1(n3090), .IN2(n3091), .IN3(n3092), .QN(n3084) );
  NAND2X0 U4599 ( .IN1(n3102), .IN2(n3114), .QN(n2629) );
  NAND3X0 U4600 ( .IN1(n3115), .IN2(n3116), .IN3(n3117), .QN(n3114) );
  AO221X1 U4601 ( .IN1(n3118), .IN2(n3121), .IN3(n3120), .IN4(n1659), .IN5(
        n3119), .Q(n3115) );
  NAND3X0 U4602 ( .IN1(n3122), .IN2(n3123), .IN3(n3124), .QN(n3116) );
  NAND2X0 U4603 ( .IN1(n3130), .IN2(n3142), .QN(n2649) );
  NAND3X0 U4604 ( .IN1(n3143), .IN2(n3144), .IN3(n3145), .QN(n3142) );
  AO221X1 U4605 ( .IN1(n3146), .IN2(n3149), .IN3(n3148), .IN4(n1678), .IN5(
        n3147), .Q(n3143) );
  NAND3X0 U4606 ( .IN1(n3150), .IN2(n3151), .IN3(n3152), .QN(n3144) );
  NAND2X0 U4607 ( .IN1(n3038), .IN2(n3039), .QN(n2794) );
  NAND3X0 U4608 ( .IN1(n3040), .IN2(n3041), .IN3(n3042), .QN(n3039) );
  AO221X1 U4609 ( .IN1(n3044), .IN2(n3047), .IN3(n3043), .IN4(n3046), .IN5(
        n3045), .Q(n3040) );
  AO221X1 U4610 ( .IN1(n3043), .IN2(n3044), .IN3(n3045), .IN4(n3046), .IN5(
        n3047), .Q(n3042) );
  NAND2X0 U4611 ( .IN1(n3070), .IN2(n3071), .QN(n2613) );
  NAND3X0 U4612 ( .IN1(n3072), .IN2(n3073), .IN3(n3074), .QN(n3071) );
  AO221X1 U4613 ( .IN1(n3076), .IN2(n3079), .IN3(n3075), .IN4(n3078), .IN5(
        n3077), .Q(n3072) );
  AO221X1 U4614 ( .IN1(n3075), .IN2(n3076), .IN3(n3077), .IN4(n3078), .IN5(
        n3079), .Q(n3074) );
  NAND2X0 U4615 ( .IN1(n3102), .IN2(n3103), .QN(n2634) );
  NAND3X0 U4616 ( .IN1(n3104), .IN2(n3105), .IN3(n3106), .QN(n3103) );
  AO221X1 U4617 ( .IN1(n3108), .IN2(n3111), .IN3(n3107), .IN4(n3110), .IN5(
        n3109), .Q(n3104) );
  AO221X1 U4618 ( .IN1(n3107), .IN2(n3108), .IN3(n3109), .IN4(n3110), .IN5(
        n3111), .Q(n3106) );
  NAND2X0 U4619 ( .IN1(n3130), .IN2(n3131), .QN(n2654) );
  NAND3X0 U4620 ( .IN1(n3132), .IN2(n3133), .IN3(n3134), .QN(n3131) );
  AO221X1 U4621 ( .IN1(n3136), .IN2(n3139), .IN3(n3135), .IN4(n3138), .IN5(
        n3137), .Q(n3132) );
  AO221X1 U4622 ( .IN1(n3135), .IN2(n3136), .IN3(n3137), .IN4(n3138), .IN5(
        n3139), .Q(n3134) );
  NAND2X0 U4623 ( .IN1(n3045), .IN2(n3044), .QN(n3048) );
  NAND2X0 U4624 ( .IN1(n3077), .IN2(n3076), .QN(n3080) );
  NAND2X0 U4625 ( .IN1(n3109), .IN2(n3108), .QN(n3112) );
  NAND2X0 U4626 ( .IN1(n3137), .IN2(n3136), .QN(n3140) );
  AND3X1 U4627 ( .IN1(n2745), .IN2(n2941), .IN3(n2692), .Q(n2855) );
  XOR2X1 U4628 ( .IN1(n2743), .IN2(n2754), .Q(n2941) );
  AND3X1 U4629 ( .IN1(n2942), .IN2(n2757), .IN3(n2756), .Q(n2692) );
  XOR2X1 U4630 ( .IN1(n2564), .IN2(n2754), .Q(n2942) );
  AND3X1 U4631 ( .IN1(n2883), .IN2(n2940), .IN3(n2855), .Q(n2766) );
  XOR2X1 U4632 ( .IN1(n2556), .IN2(n2754), .Q(n2940) );
  AND4X1 U4633 ( .IN1(n3518), .IN2(n3519), .IN3(n3520), .IN4(n3521), .Q(n3505)
         );
  NAND2X0 U4634 ( .IN1(n3509), .IN2(n2132), .QN(n3518) );
  NAND3X0 U4635 ( .IN1(n3275), .IN2(n4737), .IN3(n2128), .QN(n3519) );
  NAND3X0 U4636 ( .IN1(n2131), .IN2(n4737), .IN3(n2132), .QN(n3521) );
  AND4X1 U4637 ( .IN1(n3562), .IN2(n3563), .IN3(n3564), .IN4(n3565), .Q(n3524)
         );
  NAND2X0 U4638 ( .IN1(n3539), .IN2(n2105), .QN(n3562) );
  NAND4X0 U4639 ( .IN1(n3566), .IN2(n3542), .IN3(n3567), .IN4(n4735), .QN(
        n3563) );
  NAND3X0 U4640 ( .IN1(n2104), .IN2(n4737), .IN3(n2105), .QN(n3565) );
  AND4X1 U4641 ( .IN1(n3544), .IN2(n3545), .IN3(n3546), .IN4(n3547), .Q(n3515)
         );
  NAND2X0 U4642 ( .IN1(n3526), .IN2(n2030), .QN(n3544) );
  NAND3X0 U4643 ( .IN1(n3316), .IN2(n4737), .IN3(n2026), .QN(n3545) );
  NAND3X0 U4644 ( .IN1(n2029), .IN2(n4737), .IN3(n2030), .QN(n3547) );
  AND4X1 U4645 ( .IN1(n3598), .IN2(n3599), .IN3(n3600), .IN4(n3601), .Q(n3550)
         );
  NAND2X0 U4646 ( .IN1(n3574), .IN2(n2003), .QN(n3598) );
  NAND4X0 U4647 ( .IN1(n3602), .IN2(n3577), .IN3(n3603), .IN4(n4735), .QN(
        n3599) );
  NAND3X0 U4648 ( .IN1(n2002), .IN2(n4736), .IN3(n2003), .QN(n3601) );
  AND4X1 U4649 ( .IN1(n3579), .IN2(n3580), .IN3(n3581), .IN4(n3582), .Q(n3532)
         );
  NAND2X0 U4650 ( .IN1(n3552), .IN2(n1928), .QN(n3579) );
  NAND3X0 U4651 ( .IN1(n3356), .IN2(n4736), .IN3(n1924), .QN(n3580) );
  NAND3X0 U4652 ( .IN1(n1927), .IN2(n4737), .IN3(n1928), .QN(n3582) );
  AND4X1 U4653 ( .IN1(n3632), .IN2(n3633), .IN3(n3634), .IN4(n3635), .Q(n3585)
         );
  NAND2X0 U4654 ( .IN1(n3610), .IN2(n1901), .QN(n3632) );
  NAND4X0 U4655 ( .IN1(n3636), .IN2(n3613), .IN3(n3637), .IN4(n4735), .QN(
        n3633) );
  NAND3X0 U4656 ( .IN1(n1900), .IN2(n4736), .IN3(n1901), .QN(n3635) );
  AND4X1 U4657 ( .IN1(n3615), .IN2(n3616), .IN3(n3617), .IN4(n3618), .Q(n3558)
         );
  NAND2X0 U4658 ( .IN1(n3587), .IN2(n1826), .QN(n3615) );
  NAND3X0 U4659 ( .IN1(n3395), .IN2(n4737), .IN3(n1822), .QN(n3616) );
  NAND3X0 U4660 ( .IN1(n1825), .IN2(n4736), .IN3(n1826), .QN(n3618) );
  AND4X1 U4661 ( .IN1(n3659), .IN2(n3660), .IN3(n3661), .IN4(n3662), .Q(n3621)
         );
  NAND2X0 U4662 ( .IN1(n3644), .IN2(n1797), .QN(n3659) );
  NAND4X0 U4663 ( .IN1(n3663), .IN2(n3647), .IN3(n3664), .IN4(n4735), .QN(
        n3660) );
  NAND3X0 U4664 ( .IN1(n1796), .IN2(n4736), .IN3(n1797), .QN(n3662) );
  AO221X1 U4665 ( .IN1(n2688), .IN2(n1877), .IN3(n2763), .IN4(n2690), .IN5(
        n2691), .Q(n2746) );
  XNOR2X1 U4666 ( .IN1(n2553), .IN2(n2700), .Q(n2763) );
  AND3X1 U4667 ( .IN1(n2764), .IN2(n2765), .IN3(n2766), .Q(n2700) );
  XOR2X1 U4668 ( .IN1(n2555), .IN2(n2754), .Q(n2765) );
  NAND3X0 U4669 ( .IN1(n2100), .IN2(n2098), .IN3(n2778), .QN(n2968) );
  NAND3X0 U4670 ( .IN1(n1998), .IN2(n1996), .IN3(n2597), .QN(n2972) );
  NAND3X0 U4671 ( .IN1(n1896), .IN2(n1894), .IN3(n2618), .QN(n2976) );
  NAND3X0 U4672 ( .IN1(n1792), .IN2(n1790), .IN3(n2638), .QN(n2979) );
  AND4X1 U4673 ( .IN1(n1565), .IN2(n2235), .IN3(n2236), .IN4(n2237), .Q(n2198)
         );
  NAND2X0 U4674 ( .IN1(n2238), .IN2(n4655), .QN(n2236) );
  NAND2X0 U4675 ( .IN1(n2215), .IN2(n1956), .QN(n2235) );
  AND4X1 U4676 ( .IN1(n1565), .IN2(n2205), .IN3(n2206), .IN4(n2207), .Q(n2195)
         );
  NAND2X0 U4677 ( .IN1(n2208), .IN2(n4656), .QN(n2206) );
  NAND2X0 U4678 ( .IN1(n2210), .IN2(n1952), .QN(n2205) );
  OA222X1 U4679 ( .IN1(n3279), .IN2(n3277), .IN3(n3290), .IN4(n3276), .IN5(
        n2132), .IN6(n3282), .Q(n3292) );
  OA222X1 U4680 ( .IN1(n3320), .IN2(n3318), .IN3(n3331), .IN4(n3317), .IN5(
        n2030), .IN6(n3323), .Q(n3333) );
  OA222X1 U4681 ( .IN1(n3360), .IN2(n3358), .IN3(n3371), .IN4(n3357), .IN5(
        n1928), .IN6(n3363), .Q(n3373) );
  OA222X1 U4682 ( .IN1(n3399), .IN2(n3397), .IN3(n3410), .IN4(n3396), .IN5(
        n1826), .IN6(n3402), .Q(n3412) );
  NAND4X0 U4683 ( .IN1(n3043), .IN2(n1697), .IN3(n1702), .IN4(n3061), .QN(
        n2827) );
  INVX0 U4684 ( .IN(n3048), .QN(n1702) );
  NOR3X0 U4685 ( .IN1(n3058), .IN2(n3049), .IN3(n3059), .QN(n3061) );
  NAND4X0 U4686 ( .IN1(n3075), .IN2(n1640), .IN3(n1645), .IN4(n3093), .QN(
        n2837) );
  INVX0 U4687 ( .IN(n3080), .QN(n1645) );
  NOR3X0 U4688 ( .IN1(n3090), .IN2(n3081), .IN3(n3091), .QN(n3093) );
  NAND4X0 U4689 ( .IN1(n3107), .IN2(n1659), .IN3(n1664), .IN4(n3125), .QN(
        n2807) );
  INVX0 U4690 ( .IN(n3112), .QN(n1664) );
  NOR3X0 U4691 ( .IN1(n3122), .IN2(n3113), .IN3(n3123), .QN(n3125) );
  NAND3X0 U4692 ( .IN1(n3270), .IN2(n3277), .IN3(n3279), .QN(n3282) );
  NAND3X0 U4693 ( .IN1(n3311), .IN2(n3318), .IN3(n3320), .QN(n3323) );
  NAND3X0 U4694 ( .IN1(n3351), .IN2(n3358), .IN3(n3360), .QN(n3363) );
  NAND3X0 U4695 ( .IN1(n3390), .IN2(n3397), .IN3(n3399), .QN(n3402) );
  NAND4X0 U4696 ( .IN1(n2900), .IN2(n2708), .IN3(n4529), .IN4(n2901), .QN(
        n2893) );
  NOR4X0 U4697 ( .IN1(n2080), .IN2(n2079), .IN3(n2076), .IN4(n2499), .QN(n2901) );
  NAND4X0 U4698 ( .IN1(n2918), .IN2(n2727), .IN3(n4530), .IN4(n2919), .QN(
        n2911) );
  NOR4X0 U4699 ( .IN1(n1978), .IN2(n1977), .IN3(n1974), .IN4(n2526), .QN(n2919) );
  NAND4X0 U4700 ( .IN1(n2936), .IN2(n2743), .IN3(n1889), .IN4(n2937), .QN(
        n2929) );
  NOR4X0 U4701 ( .IN1(n2553), .IN2(n1876), .IN3(n1873), .IN4(n2552), .QN(n2937) );
  NAND4X0 U4702 ( .IN1(n2953), .IN2(n2759), .IN3(n1785), .IN4(n2954), .QN(
        n2946) );
  NOR4X0 U4703 ( .IN1(n1772), .IN2(n1771), .IN3(n1768), .IN4(n2578), .QN(n2954) );
  AND3X1 U4704 ( .IN1(n3261), .IN2(n3262), .IN3(n3263), .Q(n3255) );
  OA22X1_S38584 U4705 ( .IN1(n3264), .IN2(n3265), .IN3(n3266), .IN4(n2131), .Q(n3263)
         );
  NAND3X0 U4706 ( .IN1(n3278), .IN2(n2131), .IN3(n2118), .QN(n3262) );
  NAND3X0 U4707 ( .IN1(n3265), .IN2(n2132), .IN3(n3280), .QN(n3261) );
  XOR2X1 U4708 ( .IN1(n2501), .IN2(n4563), .Q(n3046) );
  XOR2X1 U4709 ( .IN1(n2528), .IN2(n4565), .Q(n3078) );
  XOR2X1 U4710 ( .IN1(n2554), .IN2(n4567), .Q(n3110) );
  XOR2X1 U4711 ( .IN1(n2580), .IN2(n4569), .Q(n3138) );
  XNOR2X1 U4712 ( .IN1(n2499), .IN2(n2666), .Q(n3055) );
  XNOR2X1 U4713 ( .IN1(n2526), .IN2(n2681), .Q(n3087) );
  XNOR2X1 U4714 ( .IN1(n2552), .IN2(n2696), .Q(n3119) );
  XNOR2X1 U4715 ( .IN1(n2578), .IN2(n2714), .Q(n3147) );
  XOR2X1 U4716 ( .IN1(n2553), .IN2(n1877), .Q(n3109) );
  XOR2X1 U4717 ( .IN1(n2500), .IN2(n3062), .Q(n3045) );
  XOR2X1 U4718 ( .IN1(n2527), .IN2(n3094), .Q(n3077) );
  XOR2X1 U4719 ( .IN1(n2579), .IN2(n3154), .Q(n3137) );
  INVX0 U4720 ( .IN(n4776), .QN(n4774) );
  XOR2X1 U4721 ( .IN1(n2502), .IN2(n4287), .Q(n3056) );
  XOR2X1 U4722 ( .IN1(n2529), .IN2(n4288), .Q(n3088) );
  XOR2X1 U4723 ( .IN1(n2555), .IN2(n4289), .Q(n3120) );
  XOR2X1 U4724 ( .IN1(n2581), .IN2(n4290), .Q(n3148) );
  NAND4X0 U4725 ( .IN1(n2076), .IN2(n2078), .IN3(n2499), .IN4(n2902), .QN(
        n2489) );
  AND3X1 U4726 ( .IN1(n2900), .IN2(n2079), .IN3(n2080), .Q(n2902) );
  NAND4X0 U4727 ( .IN1(n1974), .IN2(n1976), .IN3(n2526), .IN4(n2920), .QN(
        n2516) );
  AND3X1 U4728 ( .IN1(n2918), .IN2(n1977), .IN3(n1978), .Q(n2920) );
  NAND4X0 U4729 ( .IN1(n1768), .IN2(n1770), .IN3(n2578), .IN4(n2955), .QN(
        n2568) );
  AND3X1 U4730 ( .IN1(n2953), .IN2(n1771), .IN3(n1772), .Q(n2955) );
  NAND4X0 U4731 ( .IN1(n1873), .IN2(n1875), .IN3(n2552), .IN4(n2938), .QN(
        n2542) );
  AND3X1 U4732 ( .IN1(n2936), .IN2(n1876), .IN3(n2553), .Q(n2938) );
  AO21X1 U4733 ( .IN1(n3036), .IN2(n3037), .IN3(n3030), .Q(n3029) );
  NAND2X0 U4734 ( .IN1(n2096), .IN2(n1687), .QN(n3036) );
  NAND3X0 U4735 ( .IN1(n2787), .IN2(n2100), .IN3(n2790), .QN(n3037) );
  AO21X1 U4736 ( .IN1(n3068), .IN2(n3069), .IN3(n3034), .Q(n3033) );
  NAND2X0 U4737 ( .IN1(n1994), .IN2(n1630), .QN(n3068) );
  NAND3X0 U4738 ( .IN1(n2606), .IN2(n1998), .IN3(n2609), .QN(n3069) );
  AO21X1 U4739 ( .IN1(n3100), .IN2(n3101), .IN3(n3066), .Q(n3065) );
  NAND2X0 U4740 ( .IN1(n1892), .IN2(n1649), .QN(n3100) );
  NAND3X0 U4741 ( .IN1(n2627), .IN2(n1896), .IN3(n2630), .QN(n3101) );
  AO21X1 U4742 ( .IN1(n3128), .IN2(n3129), .IN3(n3098), .Q(n3097) );
  NAND2X0 U4743 ( .IN1(n1788), .IN2(n1668), .QN(n3128) );
  NAND3X0 U4744 ( .IN1(n2647), .IN2(n1792), .IN3(n2650), .QN(n3129) );
  OA22X1_S38584 U4745 ( .IN1(n2132), .IN2(n3265), .IN3(n2116), .IN4(n3279), .Q(n3267)
         );
  XOR2X1 U4746 ( .IN1(n1889), .IN2(n2563), .Q(n2883) );
  XOR2X1 U4747 ( .IN1(n2754), .IN2(n2554), .Q(n2764) );
  AO221X1 U4748 ( .IN1(n3054), .IN2(n1697), .IN3(n3055), .IN4(n3056), .IN5(
        n3057), .Q(n3053) );
  AO221X1 U4749 ( .IN1(n3086), .IN2(n1640), .IN3(n3087), .IN4(n3088), .IN5(
        n3089), .Q(n3085) );
  AO221X1 U4750 ( .IN1(n3118), .IN2(n1659), .IN3(n3119), .IN4(n3120), .IN5(
        n3121), .Q(n3117) );
  AO221X1 U4751 ( .IN1(n3146), .IN2(n1678), .IN3(n3147), .IN4(n3148), .IN5(
        n3149), .Q(n3145) );
  OA21X1 U4752 ( .IN1(n2127), .IN2(n2116), .IN3(n3279), .Q(n3269) );
  NAND4X0 U4753 ( .IN1(n1567), .IN2(n2297), .IN3(n2298), .IN4(n2279), .QN(
        n2261) );
  NAND2X0 U4754 ( .IN1(n2299), .IN2(n4658), .QN(n2298) );
  NAND2X0 U4755 ( .IN1(n2282), .IN2(n2051), .QN(n2297) );
  NAND4X0 U4756 ( .IN1(n1565), .IN2(n2225), .IN3(n2226), .IN4(n2207), .QN(
        n2189) );
  NAND2X0 U4757 ( .IN1(n2227), .IN2(n4656), .QN(n2226) );
  NAND2X0 U4758 ( .IN1(n2210), .IN2(n1949), .QN(n2225) );
  NOR2X0 U4759 ( .IN1(n3859), .IN2(n4354), .QN(n4130) );
  NAND4X0 U4760 ( .IN1(n1567), .IN2(n2319), .IN3(n2320), .IN4(n2309), .QN(
        n2260) );
  NAND2X0 U4761 ( .IN1(n2321), .IN2(n4657), .QN(n2320) );
  NAND2X0 U4762 ( .IN1(n2287), .IN2(n2049), .QN(n2319) );
  NAND4X0 U4763 ( .IN1(n1565), .IN2(n2247), .IN3(n2248), .IN4(n2237), .QN(
        n2188) );
  NAND2X0 U4764 ( .IN1(n2249), .IN2(n4655), .QN(n2248) );
  NAND2X0 U4765 ( .IN1(n2215), .IN2(n1947), .QN(n2247) );
  OA21X1 U4766 ( .IN1(n2827), .IN2(n2082), .IN3(n2791), .Q(n2786) );
  OA21X1 U4767 ( .IN1(n2837), .IN2(n1980), .IN3(n2610), .Q(n2605) );
  OA21X1 U4768 ( .IN1(n2807), .IN2(n1878), .IN3(n2631), .Q(n2626) );
  OA21X1 U4769 ( .IN1(n2817), .IN2(n1774), .IN3(n2651), .Q(n2646) );
  OA22X1_S38584 U4770 ( .IN1(n2780), .IN2(n2781), .IN3(n2782), .IN4(n2100), .Q(n2779)
         );
  NOR2X0 U4771 ( .IN1(n2098), .IN2(n2095), .QN(n2782) );
  OA22X1_S38584 U4772 ( .IN1(n2599), .IN2(n2600), .IN3(n2601), .IN4(n1998), .Q(n2598)
         );
  NOR2X0 U4773 ( .IN1(n1996), .IN2(n1993), .QN(n2601) );
  OA22X1_S38584 U4774 ( .IN1(n2640), .IN2(n2641), .IN3(n2642), .IN4(n1792), .Q(n2639)
         );
  NOR2X0 U4775 ( .IN1(n1790), .IN2(n1787), .QN(n2642) );
  NAND2X0 U4776 ( .IN1(n3038), .IN2(n2827), .QN(n2795) );
  NAND2X0 U4777 ( .IN1(n3070), .IN2(n2837), .QN(n2614) );
  NAND2X0 U4778 ( .IN1(n3102), .IN2(n2807), .QN(n2635) );
  NAND2X0 U4779 ( .IN1(n3130), .IN2(n2817), .QN(n2655) );
  NAND2X0 U4780 ( .IN1(n2778), .IN2(n2828), .QN(n2824) );
  OR3X1 U4781 ( .IN1(n2829), .IN2(n2098), .IN3(n4385), .Q(n2828) );
  NAND2X0 U4782 ( .IN1(n2597), .IN2(n2838), .QN(n2834) );
  OR3X1 U4783 ( .IN1(n2839), .IN2(n1996), .IN3(n4386), .Q(n2838) );
  NAND2X0 U4784 ( .IN1(n2618), .IN2(n2808), .QN(n2804) );
  OR3X1 U4785 ( .IN1(n2809), .IN2(n1894), .IN3(n4387), .Q(n2808) );
  NAND2X0 U4786 ( .IN1(n2638), .IN2(n2818), .QN(n2814) );
  OR3X1 U4787 ( .IN1(n2819), .IN2(n1790), .IN3(n4388), .Q(n2818) );
  INVX0 U4788 ( .IN(n2787), .QN(n2098) );
  INVX0 U4789 ( .IN(n2606), .QN(n1996) );
  INVX0 U4790 ( .IN(n2627), .QN(n1894) );
  INVX0 U4791 ( .IN(n2647), .QN(n1790) );
  INVX0 U4792 ( .IN(n2618), .QN(n1891) );
  OA22X1_S38584 U4793 ( .IN1(n3267), .IN2(n3268), .IN3(n3269), .IN4(n3270), .Q(n3266)
         );
  AOI221X1 U4794 ( .IN1(n2688), .IN2(n2696), .IN3(n2690), .IN4(n2697), .IN5(
        n2698), .QN(n2678) );
  XNOR2X1 U4795 ( .IN1(n2552), .IN2(n2699), .Q(n2697) );
  NAND2X0 U4796 ( .IN1(n2700), .IN2(n2701), .QN(n2699) );
  XOR2X1 U4797 ( .IN1(n2553), .IN2(n1889), .Q(n2701) );
  AOI221X1 U4798 ( .IN1(n1688), .IN2(n4287), .IN3(n2661), .IN4(n2857), .IN5(
        n1689), .QN(n2846) );
  XOR2X1 U4799 ( .IN1(n2502), .IN2(n2858), .Q(n2857) );
  NAND2X0 U4800 ( .IN1(n2736), .IN2(n2734), .QN(n2858) );
  AOI221X1 U4801 ( .IN1(n1688), .IN2(n4555), .IN3(n2661), .IN4(n2865), .IN5(
        n1689), .QN(n2851) );
  XOR2X1 U4802 ( .IN1(n2503), .IN2(n2866), .Q(n2865) );
  NAND2X0 U4803 ( .IN1(n2843), .IN2(n2867), .QN(n2866) );
  AOI221X1 U4804 ( .IN1(n2659), .IN2(n4389), .IN3(n2661), .IN4(n2707), .IN5(
        n2668), .QN(n2680) );
  XOR2X1 U4805 ( .IN1(n2708), .IN2(n2709), .Q(n2707) );
  NAND2X0 U4806 ( .IN1(n2663), .IN2(n2710), .QN(n2709) );
  AOI221X1 U4807 ( .IN1(n2659), .IN2(n4373), .IN3(n2661), .IN4(n2721), .IN5(
        n2668), .QN(n2694) );
  XOR2X1 U4808 ( .IN1(n2512), .IN2(n2723), .Q(n2721) );
  NAND2X0 U4809 ( .IN1(n2724), .IN2(n2725), .QN(n2723) );
  AOI221X1 U4810 ( .IN1(n1631), .IN2(n4288), .IN3(n2675), .IN4(n2868), .IN5(
        n1632), .QN(n2853) );
  XOR2X1 U4811 ( .IN1(n2529), .IN2(n2869), .Q(n2868) );
  NAND2X0 U4812 ( .IN1(n2751), .IN2(n2749), .QN(n2869) );
  AOI221X1 U4813 ( .IN1(n1631), .IN2(n4557), .IN3(n2675), .IN4(n2873), .IN5(
        n1632), .QN(n2859) );
  XOR2X1 U4814 ( .IN1(n2530), .IN2(n2874), .Q(n2873) );
  NAND2X0 U4815 ( .IN1(n2848), .IN2(n2875), .QN(n2874) );
  AOI221X1 U4816 ( .IN1(n2673), .IN2(n4390), .IN3(n2675), .IN4(n2726), .IN5(
        n2683), .QN(n2695) );
  XOR2X1 U4817 ( .IN1(n2727), .IN2(n2728), .Q(n2726) );
  NAND2X0 U4818 ( .IN1(n2677), .IN2(n2729), .QN(n2728) );
  AOI221X1 U4819 ( .IN1(n2673), .IN2(n4374), .IN3(n2675), .IN4(n2737), .IN5(
        n2683), .QN(n2712) );
  XOR2X1 U4820 ( .IN1(n2538), .IN2(n2739), .Q(n2737) );
  NAND2X0 U4821 ( .IN1(n2740), .IN2(n2741), .QN(n2739) );
  AOI221X1 U4822 ( .IN1(n1650), .IN2(n4289), .IN3(n2690), .IN4(n2876), .IN5(
        n1651), .QN(n2861) );
  XOR2X1 U4823 ( .IN1(n2555), .IN2(n2877), .Q(n2876) );
  NAND2X0 U4824 ( .IN1(n2766), .IN2(n2764), .QN(n2877) );
  AOI221X1 U4825 ( .IN1(n1650), .IN2(n4559), .IN3(n2690), .IN4(n2881), .IN5(
        n1651), .QN(n2870) );
  XOR2X1 U4826 ( .IN1(n2556), .IN2(n2882), .Q(n2881) );
  NAND2X0 U4827 ( .IN1(n2855), .IN2(n2883), .QN(n2882) );
  AOI221X1 U4828 ( .IN1(n2688), .IN2(n4391), .IN3(n2690), .IN4(n2742), .IN5(
        n2698), .QN(n2713) );
  XOR2X1 U4829 ( .IN1(n2743), .IN2(n2744), .Q(n2742) );
  NAND2X0 U4830 ( .IN1(n2692), .IN2(n2745), .QN(n2744) );
  AOI221X1 U4831 ( .IN1(n2688), .IN2(n4375), .IN3(n2690), .IN4(n2752), .IN5(
        n2698), .QN(n2731) );
  XOR2X1 U4832 ( .IN1(n2564), .IN2(n2755), .Q(n2752) );
  NAND2X0 U4833 ( .IN1(n2756), .IN2(n2757), .QN(n2755) );
  AOI221X1 U4834 ( .IN1(n1669), .IN2(n4290), .IN3(n2704), .IN4(n2884), .IN5(
        n1670), .QN(n2872) );
  XOR2X1 U4835 ( .IN1(n2581), .IN2(n2885), .Q(n2884) );
  NAND2X0 U4836 ( .IN1(n2775), .IN2(n2773), .QN(n2885) );
  AOI221X1 U4837 ( .IN1(n1669), .IN2(n4561), .IN3(n2704), .IN4(n2887), .IN5(
        n1670), .QN(n2878) );
  XOR2X1 U4838 ( .IN1(n2582), .IN2(n2888), .Q(n2887) );
  NAND2X0 U4839 ( .IN1(n2863), .IN2(n2889), .QN(n2888) );
  AOI221X1 U4840 ( .IN1(n2702), .IN2(n4392), .IN3(n2704), .IN4(n2758), .IN5(
        n2716), .QN(n2732) );
  XOR2X1 U4841 ( .IN1(n2759), .IN2(n2760), .Q(n2758) );
  NAND2X0 U4842 ( .IN1(n2706), .IN2(n2761), .QN(n2760) );
  AOI221X1 U4843 ( .IN1(n2702), .IN2(n4376), .IN3(n2704), .IN4(n2767), .IN5(
        n2716), .QN(n2747) );
  XOR2X1 U4844 ( .IN1(n2590), .IN2(n2769), .Q(n2767) );
  NAND2X0 U4845 ( .IN1(n2770), .IN2(n2771), .QN(n2769) );
  NAND2X0 U4846 ( .IN1(n2623), .IN2(n1896), .QN(n2621) );
  NAND3X0 U4847 ( .IN1(n2624), .IN2(n2625), .IN3(n2618), .QN(n2623) );
  NAND3X0 U4848 ( .IN1(n2631), .IN2(n1894), .IN3(n2632), .QN(n2624) );
  NAND4X0 U4849 ( .IN1(n2626), .IN2(n2627), .IN3(n2628), .IN4(n2629), .QN(
        n2625) );
  OA222X1 U4850 ( .IN1(n2116), .IN2(n3284), .IN3(n3277), .IN4(n3285), .IN5(
        n3275), .IN6(n3286), .Q(n3253) );
  NAND2X0 U4851 ( .IN1(n3291), .IN2(n2132), .QN(n3285) );
  OA22X1_S38584 U4852 ( .IN1(n3271), .IN2(n3270), .IN3(n3287), .IN4(n3265), .Q(n3286)
         );
  OA22X1_S38584 U4853 ( .IN1(n3273), .IN2(n3268), .IN3(n3292), .IN4(n2131), .Q(n3284)
         );
  OA222X1 U4854 ( .IN1(n2014), .IN2(n3325), .IN3(n3318), .IN4(n3326), .IN5(
        n3316), .IN6(n3327), .Q(n3294) );
  NAND2X0 U4855 ( .IN1(n3332), .IN2(n2030), .QN(n3326) );
  OA22X1_S38584 U4856 ( .IN1(n3312), .IN2(n3311), .IN3(n3328), .IN4(n3306), .Q(n3327)
         );
  OA22X1_S38584 U4857 ( .IN1(n3314), .IN2(n3309), .IN3(n3333), .IN4(n2029), .Q(n3325)
         );
  OA222X1 U4858 ( .IN1(n1912), .IN2(n3365), .IN3(n3358), .IN4(n3366), .IN5(
        n3356), .IN6(n3367), .Q(n3335) );
  NAND2X0 U4859 ( .IN1(n3372), .IN2(n1928), .QN(n3366) );
  OA22X1_S38584 U4860 ( .IN1(n3352), .IN2(n3351), .IN3(n3368), .IN4(n3346), .Q(n3367)
         );
  OA22X1_S38584 U4861 ( .IN1(n3354), .IN2(n3349), .IN3(n3373), .IN4(n1927), .Q(n3365)
         );
  OA222X1 U4862 ( .IN1(n1808), .IN2(n3404), .IN3(n3397), .IN4(n3405), .IN5(
        n3395), .IN6(n3406), .Q(n3375) );
  NAND2X0 U4863 ( .IN1(n3411), .IN2(n1826), .QN(n3405) );
  OA22X1_S38584 U4864 ( .IN1(n3391), .IN2(n3390), .IN3(n3407), .IN4(n3385), .Q(n3406)
         );
  OA22X1_S38584 U4865 ( .IN1(n3393), .IN2(n3388), .IN3(n3412), .IN4(n1825), .Q(n3404)
         );
  INVX0 U4866 ( .IN(n4116), .QN(n2100) );
  INVX0 U4867 ( .IN(n4117), .QN(n1998) );
  INVX0 U4868 ( .IN(n4118), .QN(n1896) );
  INVX0 U4869 ( .IN(n4119), .QN(n1792) );
  NAND3X0 U4870 ( .IN1(n3874), .IN2(n3875), .IN3(n3876), .QN(n3867) );
  XOR2X1 U4871 ( .IN1(n4319), .IN2(n3879), .Q(n3874) );
  XOR2X1 U4872 ( .IN1(n4377), .IN2(n3878), .Q(n3875) );
  XOR2X1 U4873 ( .IN1(n4373), .IN2(n3877), .Q(n3876) );
  NAND3X0 U4874 ( .IN1(n3771), .IN2(n3772), .IN3(n3773), .QN(n3764) );
  XOR2X1 U4875 ( .IN1(n4320), .IN2(n3776), .Q(n3771) );
  XOR2X1 U4876 ( .IN1(n4378), .IN2(n3775), .Q(n3772) );
  XOR2X1 U4877 ( .IN1(n4374), .IN2(n3774), .Q(n3773) );
  NAND3X0 U4878 ( .IN1(n3801), .IN2(n3802), .IN3(n3803), .QN(n3794) );
  XOR2X1 U4879 ( .IN1(n4321), .IN2(n3806), .Q(n3801) );
  XOR2X1 U4880 ( .IN1(n4379), .IN2(n3805), .Q(n3802) );
  XOR2X1 U4881 ( .IN1(n4375), .IN2(n3804), .Q(n3803) );
  NAND3X0 U4882 ( .IN1(n3829), .IN2(n3830), .IN3(n3831), .QN(n3822) );
  XOR2X1 U4883 ( .IN1(n4322), .IN2(n3834), .Q(n3829) );
  XOR2X1 U4884 ( .IN1(n4380), .IN2(n3833), .Q(n3830) );
  XOR2X1 U4885 ( .IN1(n4376), .IN2(n3832), .Q(n3831) );
  NAND3X0 U4886 ( .IN1(n2787), .IN2(n2095), .IN3(n2786), .QN(n2825) );
  NAND3X0 U4887 ( .IN1(n2606), .IN2(n1993), .IN3(n2605), .QN(n2835) );
  NAND3X0 U4888 ( .IN1(n2627), .IN2(n1891), .IN3(n2626), .QN(n2805) );
  NAND3X0 U4889 ( .IN1(n2647), .IN2(n1787), .IN3(n2646), .QN(n2815) );
  AOI221X1 U4890 ( .IN1(n2213), .IN2(n4655), .IN3(n2215), .IN4(n1954), .IN5(
        n2216), .QN(n2193) );
  NAND3X0 U4891 ( .IN1(n3048), .IN2(n3049), .IN3(n1699), .QN(n3041) );
  INVX0 U4892 ( .IN(n3043), .QN(n1699) );
  NAND3X0 U4893 ( .IN1(n3080), .IN2(n3081), .IN3(n1642), .QN(n3073) );
  INVX0 U4894 ( .IN(n3075), .QN(n1642) );
  NAND3X0 U4895 ( .IN1(n3112), .IN2(n3113), .IN3(n1661), .QN(n3105) );
  INVX0 U4896 ( .IN(n3107), .QN(n1661) );
  NAND3X0 U4897 ( .IN1(n3140), .IN2(n3141), .IN3(n1680), .QN(n3133) );
  INVX0 U4898 ( .IN(n3135), .QN(n1680) );
  AOI221X1 U4899 ( .IN1(n2233), .IN2(n4656), .IN3(n2210), .IN4(n1948), .IN5(
        n2216), .QN(n2200) );
  NAND2X0 U4900 ( .IN1(n2822), .IN2(n2823), .QN(n2821) );
  NAND4X0 U4901 ( .IN1(n2824), .IN2(n2825), .IN3(n2826), .IN4(n2100), .QN(
        n2822) );
  NAND2X0 U4902 ( .IN1(n2832), .IN2(n2833), .QN(n2831) );
  NAND4X0 U4903 ( .IN1(n2834), .IN2(n2835), .IN3(n2836), .IN4(n1998), .QN(
        n2832) );
  ISOLANDX1 U4904 ( .D(n2800), .ISO(n2617), .Q(n2798) );
  XOR2X1 U4905 ( .IN1(n2801), .IN2(n2627), .Q(n2800) );
  NAND2X0 U4906 ( .IN1(n2802), .IN2(n2803), .QN(n2801) );
  NAND4X0 U4907 ( .IN1(n2804), .IN2(n2805), .IN3(n2806), .IN4(n1896), .QN(
        n2802) );
  NAND2X0 U4908 ( .IN1(n2812), .IN2(n2813), .QN(n2811) );
  NAND4X0 U4909 ( .IN1(n2814), .IN2(n2815), .IN3(n2816), .IN4(n1792), .QN(
        n2812) );
  NAND2X0 U4910 ( .IN1(n3056), .IN2(n3057), .QN(n3059) );
  NAND2X0 U4911 ( .IN1(n3088), .IN2(n3089), .QN(n3091) );
  NAND2X0 U4912 ( .IN1(n3120), .IN2(n3121), .QN(n3123) );
  NAND2X0 U4913 ( .IN1(n3148), .IN2(n3149), .QN(n3151) );
  AOI221X1 U4914 ( .IN1(n2895), .IN2(n2096), .IN3(n2896), .IN4(n2100), .IN5(
        n2777), .QN(n2892) );
  NOR2X0 U4915 ( .IN1(n2898), .IN2(n2899), .QN(n2895) );
  NAND2X0 U4916 ( .IN1(n2791), .IN2(n2897), .QN(n2896) );
  NAND3X0 U4917 ( .IN1(n2778), .IN2(n2107), .IN3(n2790), .QN(n2897) );
  AOI221X1 U4918 ( .IN1(n2913), .IN2(n1994), .IN3(n2914), .IN4(n1998), .IN5(
        n2596), .QN(n2910) );
  NOR2X0 U4919 ( .IN1(n2916), .IN2(n2917), .QN(n2913) );
  NAND2X0 U4920 ( .IN1(n2610), .IN2(n2915), .QN(n2914) );
  NAND3X0 U4921 ( .IN1(n2597), .IN2(n2005), .IN3(n2609), .QN(n2915) );
  AOI221X1 U4922 ( .IN1(n2931), .IN2(n1892), .IN3(n2932), .IN4(n1896), .IN5(
        n2617), .QN(n2928) );
  NOR2X0 U4923 ( .IN1(n2934), .IN2(n2935), .QN(n2931) );
  NAND2X0 U4924 ( .IN1(n2631), .IN2(n2933), .QN(n2932) );
  NAND3X0 U4925 ( .IN1(n2618), .IN2(n1903), .IN3(n2630), .QN(n2933) );
  AOI221X1 U4926 ( .IN1(n2948), .IN2(n1788), .IN3(n2949), .IN4(n1792), .IN5(
        n2637), .QN(n2945) );
  NOR2X0 U4927 ( .IN1(n2951), .IN2(n2952), .QN(n2948) );
  NAND2X0 U4928 ( .IN1(n2651), .IN2(n2950), .QN(n2949) );
  NAND3X0 U4929 ( .IN1(n2638), .IN2(n1799), .IN3(n2650), .QN(n2950) );
  ISOLANDX1 U4930 ( .D(n2616), .ISO(n2617), .Q(n2594) );
  XOR2X1 U4931 ( .IN1(n2618), .IN2(n2619), .Q(n2616) );
  OA22X1_S38584 U4932 ( .IN1(n2620), .IN2(n2621), .IN3(n2622), .IN4(n1896), .Q(n2619)
         );
  NOR2X0 U4933 ( .IN1(n1894), .IN2(n1891), .QN(n2622) );
  NAND2X0 U4934 ( .IN1(n3047), .IN2(n3046), .QN(n3049) );
  NAND2X0 U4935 ( .IN1(n3079), .IN2(n3078), .QN(n3081) );
  NAND2X0 U4936 ( .IN1(n3111), .IN2(n3110), .QN(n3113) );
  NAND2X0 U4937 ( .IN1(n3139), .IN2(n3138), .QN(n3141) );
  NAND2X0 U4938 ( .IN1(n3055), .IN2(n3054), .QN(n3058) );
  NAND2X0 U4939 ( .IN1(n3087), .IN2(n3086), .QN(n3090) );
  NAND2X0 U4940 ( .IN1(n3119), .IN2(n3118), .QN(n3122) );
  NAND2X0 U4941 ( .IN1(n3147), .IN2(n3146), .QN(n3150) );
  NAND4X0 U4942 ( .IN1(n3135), .IN2(n1678), .IN3(n1683), .IN4(n3153), .QN(
        n2817) );
  INVX0 U4943 ( .IN(n3140), .QN(n1683) );
  NOR3X0 U4944 ( .IN1(n3150), .IN2(n3141), .IN3(n3151), .QN(n3153) );
  INVX0 U4945 ( .IN(n3062), .QN(n2081) );
  INVX0 U4946 ( .IN(n3094), .QN(n1979) );
  INVX0 U4947 ( .IN(n3154), .QN(n1773) );
  INVX0 U4948 ( .IN(n3227), .QN(n1877) );
  INVX0 U4949 ( .IN(n2898), .QN(n2107) );
  INVX0 U4950 ( .IN(n2916), .QN(n2005) );
  INVX0 U4951 ( .IN(n2934), .QN(n1903) );
  INVX0 U4952 ( .IN(n2951), .QN(n1799) );
  INVX0 U4953 ( .IN(n2565), .QN(n1874) );
  INVX0 U4954 ( .IN(n2551), .QN(n1876) );
  INVX0 U4955 ( .IN(n2708), .QN(n2078) );
  INVX0 U4956 ( .IN(n2727), .QN(n1976) );
  INVX0 U4957 ( .IN(n2743), .QN(n1875) );
  INVX0 U4958 ( .IN(n2759), .QN(n1770) );
  INVX0 U4959 ( .IN(n2512), .QN(n2076) );
  INVX0 U4960 ( .IN(n2538), .QN(n1974) );
  INVX0 U4961 ( .IN(n2564), .QN(n1873) );
  INVX0 U4962 ( .IN(n2590), .QN(n1768) );
  INVX0 U4963 ( .IN(n2500), .QN(n2080) );
  INVX0 U4964 ( .IN(n2527), .QN(n1978) );
  INVX0 U4965 ( .IN(n2579), .QN(n1772) );
  NOR4X0 U4966 ( .IN1(n2501), .IN2(n2503), .IN3(n2903), .IN4(n2502), .QN(n2900) );
  NAND2X0 U4967 ( .IN1(n2511), .IN2(n2077), .QN(n2903) );
  NOR4X0 U4968 ( .IN1(n2528), .IN2(n2530), .IN3(n2921), .IN4(n2529), .QN(n2918) );
  NAND2X0 U4969 ( .IN1(n2537), .IN2(n1975), .QN(n2921) );
  NOR4X0 U4970 ( .IN1(n2580), .IN2(n2582), .IN3(n2956), .IN4(n2581), .QN(n2953) );
  NAND2X0 U4971 ( .IN1(n2589), .IN2(n4513), .QN(n2956) );
  NOR4X0 U4972 ( .IN1(n2554), .IN2(n2556), .IN3(n2939), .IN4(n2555), .QN(n2936) );
  NAND2X0 U4973 ( .IN1(n2563), .IN2(n1874), .QN(n2939) );
  NAND2X0 U4974 ( .IN1(n2783), .IN2(n2100), .QN(n2781) );
  NAND3X0 U4975 ( .IN1(n2784), .IN2(n2785), .IN3(n2778), .QN(n2783) );
  NAND3X0 U4976 ( .IN1(n2791), .IN2(n2098), .IN3(n2792), .QN(n2784) );
  NAND4X0 U4977 ( .IN1(n2786), .IN2(n2787), .IN3(n2788), .IN4(n2789), .QN(
        n2785) );
  NAND2X0 U4978 ( .IN1(n2602), .IN2(n1998), .QN(n2600) );
  NAND3X0 U4979 ( .IN1(n2603), .IN2(n2604), .IN3(n2597), .QN(n2602) );
  NAND3X0 U4980 ( .IN1(n2610), .IN2(n1996), .IN3(n2611), .QN(n2603) );
  NAND4X0 U4981 ( .IN1(n2605), .IN2(n2606), .IN3(n2607), .IN4(n2608), .QN(
        n2604) );
  NAND2X0 U4982 ( .IN1(n2643), .IN2(n1792), .QN(n2641) );
  NAND3X0 U4983 ( .IN1(n2644), .IN2(n2645), .IN3(n2638), .QN(n2643) );
  NAND3X0 U4984 ( .IN1(n2651), .IN2(n1790), .IN3(n2652), .QN(n2644) );
  NAND4X0 U4985 ( .IN1(n2646), .IN2(n2647), .IN3(n2648), .IN4(n2649), .QN(
        n2645) );
  INVX0 U4986 ( .IN(n3060), .QN(n1697) );
  INVX0 U4987 ( .IN(n3092), .QN(n1640) );
  INVX0 U4988 ( .IN(n3124), .QN(n1659) );
  INVX0 U4989 ( .IN(n3152), .QN(n1678) );
  INVX0 U4990 ( .IN(n4323), .QN(n4592) );
  INVX0 U4991 ( .IN(n4312), .QN(n4591) );
  INVX0 U4992 ( .IN(n3038), .QN(n2082) );
  INVX0 U4993 ( .IN(n3070), .QN(n1980) );
  INVX0 U4994 ( .IN(n3102), .QN(n1878) );
  INVX0 U4995 ( .IN(n3130), .QN(n1774) );
  NAND4X0 U4996 ( .IN1(n3919), .IN2(n3920), .IN3(n3921), .IN4(n3922), .QN(
        g26135) );
  OA221X1 U4997 ( .IN1(n4331), .IN2(n3916), .IN3(n3917), .IN4(n4434), .IN5(
        n3926), .Q(n3919) );
  OA221X1 U4998 ( .IN1(n3907), .IN2(n4437), .IN3(n3908), .IN4(n4334), .IN5(
        n3924), .Q(n3921) );
  OA221X1 U4999 ( .IN1(n3906), .IN2(n4438), .IN3(n3905), .IN4(n4335), .IN5(
        n3923), .Q(n3922) );
  NAND4X0 U5000 ( .IN1(n3927), .IN2(n3928), .IN3(n3929), .IN4(n3930), .QN(
        g26104) );
  OA221X1 U5001 ( .IN1(n4302), .IN2(n3916), .IN3(n3917), .IN4(n4435), .IN5(
        n3943), .Q(n3927) );
  OA221X1 U5002 ( .IN1(n3907), .IN2(n4439), .IN3(n3908), .IN4(n4336), .IN5(
        n3937), .Q(n3929) );
  OA221X1 U5003 ( .IN1(n3906), .IN2(n4440), .IN3(n3905), .IN4(n4337), .IN5(
        n3931), .Q(n3930) );
  NAND2X0 U5004 ( .IN1(n2483), .IN2(n1587), .QN(n3734) );
  NAND2X0 U5005 ( .IN1(g13110), .IN2(n4679), .QN(n4031) );
  NAND2X0 U5006 ( .IN1(g13110), .IN2(n4587), .QN(n4032) );
  NAND2X0 U5007 ( .IN1(g13110), .IN2(g6837), .QN(n4034) );
  NAND2X0 U5008 ( .IN1(g13110), .IN2(n4684), .QN(n4033) );
  NAND2X0 U5009 ( .IN1(g13110), .IN2(n4589), .QN(n4037) );
  NAND2X0 U5010 ( .IN1(g13110), .IN2(g6573), .QN(n4040) );
  NAND2X0 U5011 ( .IN1(g13110), .IN2(n4689), .QN(n4038) );
  NAND2X0 U5012 ( .IN1(g13110), .IN2(n4591), .QN(n4043) );
  NAND2X0 U5013 ( .IN1(g13110), .IN2(n4592), .QN(n4046) );
  NAND2X0 U5014 ( .IN1(g13110), .IN2(n4694), .QN(n4044) );
  NAND2X0 U5015 ( .IN1(g13110), .IN2(n4593), .QN(n4049) );
  NAND2X0 U5016 ( .IN1(g13110), .IN2(g6231), .QN(n4051) );
  NOR2X0 U5017 ( .IN1(n3192), .IN2(n4385), .QN(n3186) );
  NOR2X0 U5018 ( .IN1(n3208), .IN2(n4386), .QN(n3202) );
  NOR2X0 U5019 ( .IN1(n3221), .IN2(n4387), .QN(n3218) );
  NOR2X0 U5020 ( .IN1(n3233), .IN2(n4388), .QN(n3232) );
  NAND2X0 U5021 ( .IN1(n3288), .IN2(n3279), .QN(n3271) );
  NAND2X0 U5022 ( .IN1(n3329), .IN2(n3320), .QN(n3312) );
  NAND2X0 U5023 ( .IN1(n3369), .IN2(n3360), .QN(n3352) );
  NAND2X0 U5024 ( .IN1(n3408), .IN2(n3399), .QN(n3391) );
  NAND2X0 U5025 ( .IN1(n3273), .IN2(n3288), .QN(n3290) );
  NAND2X0 U5026 ( .IN1(n3314), .IN2(n3329), .QN(n3331) );
  NAND2X0 U5027 ( .IN1(n3354), .IN2(n3369), .QN(n3371) );
  NAND2X0 U5028 ( .IN1(n3393), .IN2(n3408), .QN(n3410) );
  NAND2X0 U5029 ( .IN1(n3940), .IN2(n3705), .QN(n3698) );
  NAND2X0 U5030 ( .IN1(n3666), .IN2(n4641), .QN(n3620) );
  NAND2X0 U5031 ( .IN1(n3569), .IN2(n4608), .QN(n3523) );
  NAND2X0 U5032 ( .IN1(n3605), .IN2(n4620), .QN(n3549) );
  NAND2X0 U5033 ( .IN1(n3639), .IN2(g6712), .QN(n3584) );
  NAND2X0 U5034 ( .IN1(n3569), .IN2(n4610), .QN(n3538) );
  NAND2X0 U5035 ( .IN1(n3605), .IN2(n4622), .QN(n3573) );
  NAND2X0 U5036 ( .IN1(n3639), .IN2(g5472), .QN(n3609) );
  NAND2X0 U5037 ( .IN1(n3666), .IN2(n4643), .QN(n3643) );
  NAND2X0 U5038 ( .IN1(n3569), .IN2(n4605), .QN(n3513) );
  NAND2X0 U5039 ( .IN1(n3605), .IN2(n4617), .QN(n3530) );
  NAND2X0 U5040 ( .IN1(n3639), .IN2(n4629), .QN(n3556) );
  NAND2X0 U5041 ( .IN1(n3666), .IN2(n4639), .QN(n3591) );
  NAND2X0 U5042 ( .IN1(n3942), .IN2(n3934), .QN(n3916) );
  NAND2X0 U5043 ( .IN1(n4201), .IN2(n1579), .QN(n4194) );
  NAND2X0 U5044 ( .IN1(n4212), .IN2(n1579), .QN(n4197) );
  AND4X1 U5045 ( .IN1(n3622), .IN2(n3592), .IN3(n3623), .IN4(n3564), .Q(n3568)
         );
  NAND2X0 U5046 ( .IN1(n4742), .IN2(n2102), .QN(n3622) );
  OA22X1_S38584 U5047 ( .IN1(n2102), .IN2(n3624), .IN3(n4748), .IN4(n3594), .Q(n3623)
         );
  INVX0 U5048 ( .IN(n3566), .QN(n2102) );
  AND4X1 U5049 ( .IN1(n3649), .IN2(n3626), .IN3(n3650), .IN4(n3600), .Q(n3604)
         );
  NAND2X0 U5050 ( .IN1(n4741), .IN2(n2000), .QN(n3649) );
  OA22X1_S38584 U5051 ( .IN1(n2000), .IN2(n3651), .IN3(n4749), .IN4(n3628), .Q(n3650)
         );
  INVX0 U5052 ( .IN(n3602), .QN(n2000) );
  AND4X1 U5053 ( .IN1(n3667), .IN2(n3653), .IN3(n3668), .IN4(n3634), .Q(n3638)
         );
  NAND2X0 U5054 ( .IN1(n4740), .IN2(n1898), .QN(n3667) );
  OA22X1_S38584 U5055 ( .IN1(n1898), .IN2(n3669), .IN3(n4751), .IN4(n3655), .Q(n3668)
         );
  INVX0 U5056 ( .IN(n3636), .QN(n1898) );
  AND4X1 U5057 ( .IN1(n3674), .IN2(n3671), .IN3(n3675), .IN4(n3661), .Q(n3665)
         );
  NAND2X0 U5058 ( .IN1(n4738), .IN2(n1794), .QN(n3674) );
  OA22X1_S38584 U5059 ( .IN1(n1794), .IN2(n3676), .IN3(n4752), .IN4(n3673), .Q(n3675)
         );
  INVX0 U5060 ( .IN(n3663), .QN(n1794) );
  NAND3X0 U5061 ( .IN1(n2095), .IN2(n2098), .IN3(n4116), .QN(n2504) );
  NAND3X0 U5062 ( .IN1(n1993), .IN2(n1996), .IN3(n4117), .QN(n2531) );
  NAND3X0 U5063 ( .IN1(n1891), .IN2(n1894), .IN3(n4118), .QN(n2557) );
  NAND3X0 U5064 ( .IN1(n1787), .IN2(n1790), .IN3(n4119), .QN(n2583) );
  AND3X1 U5065 ( .IN1(n3535), .IN2(n3536), .IN3(n3537), .Q(n3511) );
  NAND3X0 U5066 ( .IN1(n2129), .IN2(n4737), .IN3(n3275), .QN(n3536) );
  AND3X1 U5067 ( .IN1(n3570), .IN2(n3571), .IN3(n3572), .Q(n3528) );
  NAND3X0 U5068 ( .IN1(n2027), .IN2(n4737), .IN3(n3316), .QN(n3571) );
  AND3X1 U5069 ( .IN1(n3606), .IN2(n3607), .IN3(n3608), .Q(n3554) );
  NAND3X0 U5070 ( .IN1(n1925), .IN2(n4737), .IN3(n3356), .QN(n3607) );
  AND3X1 U5071 ( .IN1(n3653), .IN2(n3654), .IN3(n3655), .Q(n3614) );
  NAND3X0 U5072 ( .IN1(n1899), .IN2(n4737), .IN3(n3613), .QN(n3654) );
  AND3X1 U5073 ( .IN1(n3640), .IN2(n3641), .IN3(n3642), .Q(n3589) );
  NAND3X0 U5074 ( .IN1(n1823), .IN2(n4736), .IN3(n3395), .QN(n3641) );
  AND3X1 U5075 ( .IN1(n3671), .IN2(n3672), .IN3(n3673), .Q(n3648) );
  NAND3X0 U5076 ( .IN1(n1795), .IN2(n4737), .IN3(n3647), .QN(n3672) );
  OA222X1 U5077 ( .IN1(n3288), .IN2(n3276), .IN3(n2120), .IN4(n3289), .IN5(
        n3268), .IN6(n3290), .Q(n3287) );
  NAND2X0 U5078 ( .IN1(n3277), .IN2(n2129), .QN(n3289) );
  OA222X1 U5079 ( .IN1(n3329), .IN2(n3317), .IN3(n2018), .IN4(n3330), .IN5(
        n3309), .IN6(n3331), .Q(n3328) );
  NAND2X0 U5080 ( .IN1(n3318), .IN2(n2027), .QN(n3330) );
  OA222X1 U5081 ( .IN1(n3369), .IN2(n3357), .IN3(n1916), .IN4(n3370), .IN5(
        n3349), .IN6(n3371), .Q(n3368) );
  NAND2X0 U5082 ( .IN1(n3358), .IN2(n1925), .QN(n3370) );
  OA222X1 U5083 ( .IN1(n3408), .IN2(n3396), .IN3(n1812), .IN4(n3409), .IN5(
        n3388), .IN6(n3410), .Q(n3407) );
  NAND2X0 U5084 ( .IN1(n3397), .IN2(n1823), .QN(n3409) );
  NAND2X0 U5085 ( .IN1(n3276), .IN2(n3277), .QN(n3268) );
  NAND2X0 U5086 ( .IN1(n3317), .IN2(n3318), .QN(n3309) );
  NAND2X0 U5087 ( .IN1(n3357), .IN2(n3358), .QN(n3349) );
  NAND2X0 U5088 ( .IN1(n3396), .IN2(n3397), .QN(n3388) );
  NOR3X0 U5089 ( .IN1(n2666), .IN2(n3062), .IN3(n3198), .QN(n3197) );
  NOR3X0 U5090 ( .IN1(n2681), .IN2(n3094), .IN3(n3214), .QN(n3213) );
  NOR3X0 U5091 ( .IN1(n2714), .IN2(n3154), .IN3(n3239), .QN(n3238) );
  NOR3X0 U5092 ( .IN1(n2696), .IN2(n3227), .IN3(n3228), .QN(n3226) );
  INVX0 U5093 ( .IN(g27380), .QN(n1576) );
  NOR2X0 U5094 ( .IN1(n4482), .IN2(n2483), .QN(n2484) );
  NAND2X0 U5095 ( .IN1(n1693), .IN2(n4285), .QN(n3195) );
  NAND2X0 U5096 ( .IN1(n1636), .IN2(n4284), .QN(n3211) );
  NAND2X0 U5097 ( .IN1(n1655), .IN2(n4283), .QN(n3224) );
  NAND2X0 U5098 ( .IN1(n1674), .IN2(n4282), .QN(n3236) );
  AND3X1 U5099 ( .IN1(n3302), .IN2(n3303), .IN3(n3304), .Q(n3296) );
  OA22X1_S38584 U5100 ( .IN1(n3305), .IN2(n3306), .IN3(n3307), .IN4(n2029), .Q(n3304)
         );
  NAND3X0 U5101 ( .IN1(n3319), .IN2(n2029), .IN3(n2016), .QN(n3303) );
  NAND3X0 U5102 ( .IN1(n3306), .IN2(n2030), .IN3(n3321), .QN(n3302) );
  AND3X1 U5103 ( .IN1(n3342), .IN2(n3343), .IN3(n3344), .Q(n3337) );
  OA22X1_S38584 U5104 ( .IN1(n3345), .IN2(n3346), .IN3(n3347), .IN4(n1927), .Q(n3344)
         );
  NAND3X0 U5105 ( .IN1(n3359), .IN2(n1927), .IN3(n1914), .QN(n3343) );
  NAND3X0 U5106 ( .IN1(n3346), .IN2(n1928), .IN3(n3361), .QN(n3342) );
  AND3X1 U5107 ( .IN1(n3381), .IN2(n3382), .IN3(n3383), .Q(n3377) );
  OA22X1_S38584 U5108 ( .IN1(n3384), .IN2(n3385), .IN3(n3386), .IN4(n1825), .Q(n3383)
         );
  NAND3X0 U5109 ( .IN1(n3398), .IN2(n1825), .IN3(n1810), .QN(n3382) );
  NAND3X0 U5110 ( .IN1(n3385), .IN2(n1826), .IN3(n3400), .QN(n3381) );
  AO22X1 U5111 ( .IN1(n3275), .IN2(n3276), .IN3(n3279), .IN4(n2116), .Q(n3291)
         );
  AO22X1 U5112 ( .IN1(n3316), .IN2(n3317), .IN3(n3320), .IN4(n2014), .Q(n3332)
         );
  AO22X1 U5113 ( .IN1(n3356), .IN2(n3357), .IN3(n3360), .IN4(n1912), .Q(n3372)
         );
  AO22X1 U5114 ( .IN1(n3395), .IN2(n3396), .IN3(n3399), .IN4(n1808), .Q(n3411)
         );
  INVX0 U5115 ( .IN(n4776), .QN(n4772) );
  INVX0 U5116 ( .IN(n4776), .QN(n4773) );
  INVX0 U5117 ( .IN(n4770), .QN(n4775) );
  INVX0 U5118 ( .IN(n4776), .QN(n4771) );
  INVX0 U5119 ( .IN(n4351), .QN(n4728) );
  INVX0 U5120 ( .IN(n4351), .QN(n4729) );
  INVX0 U5121 ( .IN(n4726), .QN(n4724) );
  INVX0 U5122 ( .IN(n4351), .QN(n4727) );
  INVX0 U5123 ( .IN(n4725), .QN(n4699) );
  INVX0 U5124 ( .IN(n4726), .QN(n4725) );
  OA221X1 U5125 ( .IN1(n3708), .IN2(n4331), .IN3(n1626), .IN4(n4302), .IN5(
        n4405), .Q(n3707) );
  AND3X1 U5126 ( .IN1(n4061), .IN2(n2481), .IN3(n4098), .Q(g24476) );
  NAND2X0 U5127 ( .IN1(n4099), .IN2(n4349), .QN(n4098) );
  ISOLANDX1 U5128 ( .D(n3933), .ISO(n4406), .Q(n3940) );
  NAND2X0 U5129 ( .IN1(n3279), .IN2(n2132), .QN(n3537) );
  NAND2X0 U5130 ( .IN1(n3320), .IN2(n2030), .QN(n3572) );
  NAND2X0 U5131 ( .IN1(n3360), .IN2(n1928), .QN(n3608) );
  NAND2X0 U5132 ( .IN1(n3399), .IN2(n1826), .QN(n3642) );
  NOR2X0 U5133 ( .IN1(n4398), .IN2(n4186), .QN(n4185) );
  NOR2X0 U5134 ( .IN1(n4400), .IN2(n4189), .QN(n4188) );
  NOR2X0 U5135 ( .IN1(n4402), .IN2(n4192), .QN(n4191) );
  NOR2X0 U5136 ( .IN1(n4404), .IN2(n4135), .QN(n4134) );
  OA22X1_S38584 U5137 ( .IN1(n2030), .IN2(n3306), .IN3(n2014), .IN4(n3320), .Q(n3308)
         );
  OA22X1_S38584 U5138 ( .IN1(n1928), .IN2(n3346), .IN3(n1912), .IN4(n3360), .Q(n3348)
         );
  OA22X1_S38584 U5139 ( .IN1(n1826), .IN2(n3385), .IN3(n1808), .IN4(n3399), .Q(n3387)
         );
  INVX0 U5140 ( .IN(n4169), .QN(n2088) );
  ISOLANDX1 U5141 ( .D(n3939), .ISO(n4405), .Q(n3936) );
  NAND2X0 U5142 ( .IN1(n4200), .IN2(n1629), .QN(n4195) );
  NAND2X0 U5143 ( .IN1(n4200), .IN2(n1628), .QN(n4198) );
  INVX0 U5144 ( .IN(n4171), .QN(n1986) );
  INVX0 U5145 ( .IN(n4174), .QN(n1884) );
  INVX0 U5146 ( .IN(n4177), .QN(n1780) );
  OA21X1 U5147 ( .IN1(n2025), .IN2(n2014), .IN3(n3320), .Q(n3310) );
  OA21X1 U5148 ( .IN1(n1923), .IN2(n1912), .IN3(n3360), .Q(n3350) );
  OA21X1 U5149 ( .IN1(n1821), .IN2(n1808), .IN3(n3399), .Q(n3389) );
  NOR2X0 U5150 ( .IN1(n4419), .IN2(n4106), .QN(n4105) );
  NOR2X0 U5151 ( .IN1(n4420), .IN2(n4109), .QN(n4108) );
  NOR2X0 U5152 ( .IN1(n4421), .IN2(n4112), .QN(n4111) );
  NOR2X0 U5153 ( .IN1(n4422), .IN2(n4115), .QN(n4114) );
  NOR2X0 U5154 ( .IN1(n4467), .IN2(n3681), .QN(n3680) );
  NOR2X0 U5155 ( .IN1(n4397), .IN2(n3747), .QN(n3746) );
  NOR2X0 U5156 ( .IN1(n4468), .IN2(n3489), .QN(n3488) );
  NOR2X0 U5157 ( .IN1(n4399), .IN2(n3755), .QN(n3754) );
  NOR2X0 U5158 ( .IN1(n4469), .IN2(n3493), .QN(n3492) );
  NOR2X0 U5159 ( .IN1(n4401), .IN2(n3785), .QN(n3784) );
  NOR2X0 U5160 ( .IN1(n4470), .IN2(n3497), .QN(n3496) );
  NOR2X0 U5161 ( .IN1(n4403), .IN2(n3815), .QN(n3814) );
  XNOR2X1 U5162 ( .IN1(n3192), .IN2(n3193), .Q(n3180) );
  OA21X1 U5163 ( .IN1(n1692), .IN2(n2089), .IN3(n3194), .Q(n3193) );
  INVX0 U5164 ( .IN(n3185), .QN(n1692) );
  OAI221X1 U5165 ( .IN1(n3195), .IN2(n2106), .IN3(n3196), .IN4(n2106), .IN5(
        n2090), .QN(n3194) );
  XNOR2X1 U5166 ( .IN1(n3208), .IN2(n3209), .Q(n3188) );
  OA21X1 U5167 ( .IN1(n1635), .IN2(n1987), .IN3(n3210), .Q(n3209) );
  INVX0 U5168 ( .IN(n3201), .QN(n1635) );
  OAI221X1 U5169 ( .IN1(n3211), .IN2(n2004), .IN3(n3212), .IN4(n2004), .IN5(
        n1988), .QN(n3210) );
  XNOR2X1 U5170 ( .IN1(n3221), .IN2(n3222), .Q(n3204) );
  OA21X1 U5171 ( .IN1(n1654), .IN2(n1885), .IN3(n3223), .Q(n3222) );
  INVX0 U5172 ( .IN(n3217), .QN(n1654) );
  OAI221X1 U5173 ( .IN1(n3224), .IN2(n1902), .IN3(n3225), .IN4(n1902), .IN5(
        n1886), .QN(n3223) );
  XNOR2X1 U5174 ( .IN1(n3233), .IN2(n3234), .Q(n3220) );
  OA21X1 U5175 ( .IN1(n1673), .IN2(n1781), .IN3(n3235), .Q(n3234) );
  INVX0 U5176 ( .IN(n3231), .QN(n1673) );
  OAI221X1 U5177 ( .IN1(n3236), .IN2(n1798), .IN3(n3237), .IN4(n1798), .IN5(
        n1782), .QN(n3235) );
  XOR2X1 U5178 ( .IN1(n3014), .IN2(n4283), .Q(n3005) );
  NAND2X0 U5179 ( .IN1(n3015), .IN2(n3016), .QN(n3014) );
  OR4X1 U5180 ( .IN1(n2631), .IN2(n1655), .IN3(n1885), .IN4(n4283), .Q(n3016)
         );
  AO221X1 U5181 ( .IN1(n3017), .IN2(n1906), .IN3(n4283), .IN4(n3018), .IN5(
        n3019), .Q(n3015) );
  NAND3X0 U5182 ( .IN1(n1748), .IN2(n4405), .IN3(n3942), .QN(n3699) );
  INVX0 U5183 ( .IN(n3275), .QN(n2131) );
  INVX0 U5184 ( .IN(n3316), .QN(n2029) );
  INVX0 U5185 ( .IN(n3356), .QN(n1927) );
  INVX0 U5186 ( .IN(n3395), .QN(n1825) );
  AOI22X1 U5187 ( .IN1(n3509), .IN2(n2130), .IN3(n3510), .IN4(n2130), .QN(
        n3502) );
  INVX0 U5188 ( .IN(n3271), .QN(n2130) );
  NOR2X0 U5189 ( .IN1(n4745), .IN2(n3275), .QN(n3510) );
  AOI22X1 U5190 ( .IN1(n3526), .IN2(n2028), .IN3(n3527), .IN4(n2028), .QN(
        n3506) );
  INVX0 U5191 ( .IN(n3312), .QN(n2028) );
  NOR2X0 U5192 ( .IN1(n4747), .IN2(n3316), .QN(n3527) );
  AOI22X1 U5193 ( .IN1(n3552), .IN2(n1926), .IN3(n3553), .IN4(n1926), .QN(
        n3516) );
  INVX0 U5194 ( .IN(n3352), .QN(n1926) );
  NOR2X0 U5195 ( .IN1(n4748), .IN2(n3356), .QN(n3553) );
  AOI22X1 U5196 ( .IN1(n3587), .IN2(n1824), .IN3(n3588), .IN4(n1824), .QN(
        n3533) );
  INVX0 U5197 ( .IN(n3391), .QN(n1824) );
  NOR2X0 U5198 ( .IN1(n4750), .IN2(n3395), .QN(n3588) );
  AOI22X1 U5199 ( .IN1(n3539), .IN2(n3540), .IN3(n3541), .IN4(n3540), .QN(
        n3512) );
  NOR2X0 U5200 ( .IN1(n2103), .IN2(n2105), .QN(n3540) );
  NOR2X0 U5201 ( .IN1(n4746), .IN2(n3542), .QN(n3541) );
  AOI22X1 U5202 ( .IN1(n3574), .IN2(n3575), .IN3(n3576), .IN4(n3575), .QN(
        n3529) );
  NOR2X0 U5203 ( .IN1(n2001), .IN2(n2003), .QN(n3575) );
  NOR2X0 U5204 ( .IN1(n4749), .IN2(n3577), .QN(n3576) );
  AOI22X1 U5205 ( .IN1(n3610), .IN2(n3611), .IN3(n3612), .IN4(n3611), .QN(
        n3555) );
  NOR2X0 U5206 ( .IN1(n1899), .IN2(n1901), .QN(n3611) );
  NOR2X0 U5207 ( .IN1(n4751), .IN2(n3613), .QN(n3612) );
  AOI22X1 U5208 ( .IN1(n3644), .IN2(n3645), .IN3(n3646), .IN4(n3645), .QN(
        n3590) );
  NOR2X0 U5209 ( .IN1(n1795), .IN2(n1797), .QN(n3645) );
  NOR2X0 U5210 ( .IN1(n4752), .IN2(n3647), .QN(n3646) );
  NAND2X0 U5211 ( .IN1(n3932), .IN2(n3933), .QN(n3903) );
  NAND3X0 U5212 ( .IN1(n4406), .IN2(n4329), .IN3(n3936), .QN(n3917) );
  AO21X1 U5213 ( .IN1(n3004), .IN2(n2791), .IN3(n1693), .Q(n3001) );
  AO21X1 U5214 ( .IN1(n3012), .IN2(n2610), .IN3(n1636), .Q(n3009) );
  AO21X1 U5215 ( .IN1(n3020), .IN2(n2631), .IN3(n1655), .Q(n3017) );
  AO21X1 U5216 ( .IN1(n3027), .IN2(n2651), .IN3(n1674), .Q(n3024) );
  NAND3X0 U5217 ( .IN1(n3933), .IN2(n4406), .IN3(n3939), .QN(n3912) );
  NAND3X0 U5218 ( .IN1(n2791), .IN2(n2109), .IN3(n3197), .QN(n3196) );
  NAND3X0 U5219 ( .IN1(n2610), .IN2(n2008), .IN3(n3213), .QN(n3212) );
  NAND3X0 U5220 ( .IN1(n2631), .IN2(n1906), .IN3(n3226), .QN(n3225) );
  NAND3X0 U5221 ( .IN1(n2651), .IN2(n1802), .IN3(n3238), .QN(n3237) );
  NAND3X0 U5222 ( .IN1(n1748), .IN2(n4405), .IN3(n3939), .QN(n3910) );
  INVX0 U5223 ( .IN(n3288), .QN(n2132) );
  INVX0 U5224 ( .IN(n3329), .QN(n2030) );
  INVX0 U5225 ( .IN(n3369), .QN(n1928) );
  INVX0 U5226 ( .IN(n3408), .QN(n1826) );
  NAND3X0 U5227 ( .IN1(n3004), .IN2(n3185), .IN3(n2090), .QN(n3177) );
  NAND3X0 U5228 ( .IN1(n3012), .IN2(n3201), .IN3(n1988), .QN(n3182) );
  NAND3X0 U5229 ( .IN1(n3020), .IN2(n3217), .IN3(n1886), .QN(n3190) );
  NAND3X0 U5230 ( .IN1(n3027), .IN2(n3231), .IN3(n1782), .QN(n3206) );
  INVX0 U5231 ( .IN(n3279), .QN(n2129) );
  INVX0 U5232 ( .IN(n3320), .QN(n2027) );
  INVX0 U5233 ( .IN(n3360), .QN(n1925) );
  INVX0 U5234 ( .IN(n3399), .QN(n1823) );
  NAND4X0 U5235 ( .IN1(n3566), .IN2(n3567), .IN3(n4740), .IN4(n2104), .QN(
        n3564) );
  NAND4X0 U5236 ( .IN1(n3602), .IN2(n3603), .IN3(n4741), .IN4(n2002), .QN(
        n3600) );
  NAND4X0 U5237 ( .IN1(n3636), .IN2(n3637), .IN3(n4739), .IN4(n1900), .QN(
        n3634) );
  NAND4X0 U5238 ( .IN1(n3663), .IN2(n3664), .IN3(n4738), .IN4(n1796), .QN(
        n3661) );
  OA22X1_S38584 U5239 ( .IN1(n3271), .IN2(n3272), .IN3(n3273), .IN4(n3274), .Q(n3264)
         );
  NAND2X0 U5240 ( .IN1(n2119), .IN2(n3277), .QN(n3272) );
  OA21X1 U5241 ( .IN1(n3275), .IN2(n2120), .IN3(n3276), .Q(n3274) );
  OA22X1_S38584 U5242 ( .IN1(n3312), .IN2(n3313), .IN3(n3314), .IN4(n3315), .Q(n3305)
         );
  NAND2X0 U5243 ( .IN1(n2017), .IN2(n3318), .QN(n3313) );
  OA21X1 U5244 ( .IN1(n3316), .IN2(n2018), .IN3(n3317), .Q(n3315) );
  OA22X1_S38584 U5245 ( .IN1(n3352), .IN2(n3353), .IN3(n3354), .IN4(n3355), .Q(n3345)
         );
  NAND2X0 U5246 ( .IN1(n1915), .IN2(n3358), .QN(n3353) );
  OA21X1 U5247 ( .IN1(n3356), .IN2(n1916), .IN3(n3357), .Q(n3355) );
  OA22X1_S38584 U5248 ( .IN1(n3391), .IN2(n3392), .IN3(n3393), .IN4(n3394), .Q(n3384)
         );
  NAND2X0 U5249 ( .IN1(n1811), .IN2(n3397), .QN(n3392) );
  OA21X1 U5250 ( .IN1(n3395), .IN2(n1812), .IN3(n3396), .Q(n3394) );
  OA22X1_S38584 U5251 ( .IN1(n3308), .IN2(n3309), .IN3(n3310), .IN4(n3311), .Q(n3307)
         );
  OA22X1_S38584 U5252 ( .IN1(n3348), .IN2(n3349), .IN3(n3350), .IN4(n3351), .Q(n3347)
         );
  OA22X1_S38584 U5253 ( .IN1(n3387), .IN2(n3388), .IN3(n3389), .IN4(n3390), .Q(n3386)
         );
  NAND2X0 U5254 ( .IN1(n3625), .IN2(n2105), .QN(n3594) );
  NAND2X0 U5255 ( .IN1(n3652), .IN2(n2003), .QN(n3628) );
  NAND2X0 U5256 ( .IN1(n3670), .IN2(n1901), .QN(n3655) );
  NAND2X0 U5257 ( .IN1(n3677), .IN2(n1797), .QN(n3673) );
  NOR3X0 U5258 ( .IN1(n4659), .IN2(n4303), .IN3(n3843), .QN(n3841) );
  NOR3X0 U5259 ( .IN1(n4657), .IN2(n4297), .IN3(n3845), .QN(n3842) );
  NOR3X0 U5260 ( .IN1(n4655), .IN2(n4304), .IN3(n3847), .QN(n3844) );
  NOR3X0 U5261 ( .IN1(n4653), .IN2(n4310), .IN3(n3848), .QN(n3846) );
  NAND2X0 U5262 ( .IN1(n3940), .IN2(n3942), .QN(n3703) );
  NAND2X0 U5263 ( .IN1(n1747), .IN2(n3934), .QN(n3905) );
  INVX0 U5264 ( .IN(n3277), .QN(n2118) );
  INVX0 U5265 ( .IN(n3318), .QN(n2016) );
  INVX0 U5266 ( .IN(n3358), .QN(n1914) );
  INVX0 U5267 ( .IN(n3397), .QN(n1810) );
  NAND2X0 U5268 ( .IN1(n3939), .IN2(n3940), .QN(n3907) );
  AO21X1 U5269 ( .IN1(n3445), .IN2(n3446), .IN3(n4385), .Q(n3437) );
  NAND3X0 U5270 ( .IN1(n2091), .IN2(n3449), .IN3(n2110), .QN(n3445) );
  NAND3X0 U5271 ( .IN1(n3447), .IN2(n3448), .IN3(n1691), .QN(n3446) );
  AO21X1 U5272 ( .IN1(n3457), .IN2(n3458), .IN3(n4386), .Q(n3441) );
  NAND3X0 U5273 ( .IN1(n1989), .IN2(n3461), .IN3(n2007), .QN(n3457) );
  NAND3X0 U5274 ( .IN1(n3459), .IN2(n3460), .IN3(n1634), .QN(n3458) );
  AO21X1 U5275 ( .IN1(n3469), .IN2(n3470), .IN3(n4387), .Q(n3453) );
  NAND3X0 U5276 ( .IN1(n1887), .IN2(n3473), .IN3(n1905), .QN(n3469) );
  NAND3X0 U5277 ( .IN1(n3471), .IN2(n3472), .IN3(n1653), .QN(n3470) );
  AO21X1 U5278 ( .IN1(n3478), .IN2(n3479), .IN3(n4388), .Q(n3465) );
  NAND3X0 U5279 ( .IN1(n1783), .IN2(n3482), .IN3(n1801), .QN(n3478) );
  NAND3X0 U5280 ( .IN1(n3480), .IN2(n3481), .IN3(n1672), .QN(n3479) );
  NAND2X0 U5281 ( .IN1(n3939), .IN2(n3934), .QN(n3915) );
  AND3X1 U5282 ( .IN1(n3592), .IN2(n3593), .IN3(n3594), .Q(n3543) );
  NAND3X0 U5283 ( .IN1(n2103), .IN2(n4736), .IN3(n3542), .QN(n3593) );
  AND3X1 U5284 ( .IN1(n3626), .IN2(n3627), .IN3(n3628), .Q(n3578) );
  NAND3X0 U5285 ( .IN1(n2001), .IN2(n4736), .IN3(n3577), .QN(n3627) );
  INVX0 U5286 ( .IN(g25435), .QN(n1573) );
  INVX0 U5287 ( .IN(n3542), .QN(n2104) );
  INVX0 U5288 ( .IN(n3577), .QN(n2002) );
  INVX0 U5289 ( .IN(n3613), .QN(n1900) );
  INVX0 U5290 ( .IN(n3647), .QN(n1796) );
  NAND2X0 U5291 ( .IN1(n3934), .IN2(n3705), .QN(n3695) );
  INVX0 U5292 ( .IN(n4285), .QN(n2109) );
  INVX0 U5293 ( .IN(n4284), .QN(n2008) );
  INVX0 U5294 ( .IN(n4283), .QN(n1906) );
  INVX0 U5295 ( .IN(n4282), .QN(n1802) );
  NBUFFX2 U5296 ( .IN(n2353), .Q(n4660) );
  NBUFFX2 U5297 ( .IN(n2281), .Q(n4658) );
  NBUFFX2 U5298 ( .IN(n2209), .Q(n4656) );
  NBUFFX2 U5299 ( .IN(n2432), .Q(n4654) );
  INVX0 U5300 ( .IN(n2365), .QN(n2137) );
  INVX0 U5301 ( .IN(n2293), .QN(n2035) );
  INVX0 U5302 ( .IN(n2221), .QN(n1933) );
  INVX0 U5303 ( .IN(n2455), .QN(n1833) );
  NBUFFX2 U5304 ( .IN(n2358), .Q(n4659) );
  NBUFFX2 U5305 ( .IN(n2286), .Q(n4657) );
  NBUFFX2 U5306 ( .IN(n2214), .Q(n4655) );
  NBUFFX2 U5307 ( .IN(n2437), .Q(n4653) );
  OR2X1 U5308 ( .IN1(n4099), .IN2(n4349), .Q(n4061) );
  INVX0 U5309 ( .IN(n3567), .QN(n2105) );
  INVX0 U5310 ( .IN(n3603), .QN(n2003) );
  INVX0 U5311 ( .IN(n3637), .QN(n1901) );
  INVX0 U5312 ( .IN(n3664), .QN(n1797) );
  INVX0 U5313 ( .IN(n3276), .QN(n2119) );
  INVX0 U5314 ( .IN(n3317), .QN(n2017) );
  INVX0 U5315 ( .IN(n3357), .QN(n1915) );
  INVX0 U5316 ( .IN(n3396), .QN(n1811) );
  INVX0 U5317 ( .IN(g24734), .QN(n1572) );
  XOR2X1 U5318 ( .IN1(n4397), .IN2(n2158), .Q(n3961) );
  XOR2X1 U5319 ( .IN1(n4399), .IN2(n2056), .Q(n3981) );
  XOR2X1 U5320 ( .IN1(n4401), .IN2(n1954), .Q(n4003) );
  XOR2X1 U5321 ( .IN1(n4403), .IN2(n1853), .Q(n4021) );
  XOR2X1 U5322 ( .IN1(n4398), .IN2(n2157), .Q(n3960) );
  XOR2X1 U5323 ( .IN1(n4400), .IN2(n2055), .Q(n3980) );
  XOR2X1 U5324 ( .IN1(n4402), .IN2(n1953), .Q(n4002) );
  XOR2X1 U5325 ( .IN1(n4404), .IN2(n1852), .Q(n4020) );
  XOR2X1 U5326 ( .IN1(n4408), .IN2(n2156), .Q(n3959) );
  XOR2X1 U5327 ( .IN1(n4410), .IN2(n2054), .Q(n3979) );
  XOR2X1 U5328 ( .IN1(n4412), .IN2(n1952), .Q(n4001) );
  XOR2X1 U5329 ( .IN1(n4414), .IN2(n1851), .Q(n4019) );
  INVX0 U5330 ( .IN(n3314), .QN(n2025) );
  INVX0 U5331 ( .IN(n3354), .QN(n1923) );
  INVX0 U5332 ( .IN(n3393), .QN(n1821) );
  INVX0 U5333 ( .IN(n3273), .QN(n2127) );
  NAND2X0 U5334 ( .IN1(n2481), .IN2(n2482), .QN(n4273) );
  AO21X1 U5335 ( .IN1(n4482), .IN2(n2483), .IN3(n2484), .Q(n2482) );
  XOR2X1 U5336 ( .IN1(n2419), .IN2(n2420), .Q(n4260) );
  XOR2X1 U5337 ( .IN1(n2419), .IN2(n2421), .Q(n4261) );
  INVX0 U5338 ( .IN(n3448), .QN(n2110) );
  INVX0 U5339 ( .IN(n3460), .QN(n2007) );
  INVX0 U5340 ( .IN(n3472), .QN(n1905) );
  INVX0 U5341 ( .IN(n3481), .QN(n1801) );
  INVX0 U5342 ( .IN(n3265), .QN(n2116) );
  INVX0 U5343 ( .IN(n3306), .QN(n2014) );
  INVX0 U5344 ( .IN(n3346), .QN(n1912) );
  INVX0 U5345 ( .IN(n3385), .QN(n1808) );
  NAND4X0 U5346 ( .IN1(n3965), .IN2(n3966), .IN3(n3967), .IN4(n3968), .QN(
        n3957) );
  XOR2X1 U5347 ( .IN1(n4407), .IN2(n2152), .Q(n3966) );
  XOR2X1 U5348 ( .IN1(n4393), .IN2(n2151), .Q(n3965) );
  XOR2X1 U5349 ( .IN1(n4415), .IN2(n2153), .Q(n3967) );
  NAND4X0 U5350 ( .IN1(n3985), .IN2(n3986), .IN3(n3987), .IN4(n3988), .QN(
        n3977) );
  XOR2X1 U5351 ( .IN1(n4409), .IN2(n2050), .Q(n3986) );
  XOR2X1 U5352 ( .IN1(n4394), .IN2(n2049), .Q(n3985) );
  XOR2X1 U5353 ( .IN1(n4416), .IN2(n2051), .Q(n3987) );
  NAND4X0 U5354 ( .IN1(n4007), .IN2(n4008), .IN3(n4009), .IN4(n4010), .QN(
        n3999) );
  XOR2X1 U5355 ( .IN1(n4411), .IN2(n1948), .Q(n4008) );
  XOR2X1 U5356 ( .IN1(n4395), .IN2(n1947), .Q(n4007) );
  XOR2X1 U5357 ( .IN1(n4417), .IN2(n1949), .Q(n4009) );
  NAND4X0 U5358 ( .IN1(n4025), .IN2(n4026), .IN3(n4027), .IN4(n4028), .QN(
        n4017) );
  XOR2X1 U5359 ( .IN1(n4413), .IN2(n1847), .Q(n4026) );
  XOR2X1 U5360 ( .IN1(n4396), .IN2(n1846), .Q(n4025) );
  XOR2X1 U5361 ( .IN1(n4418), .IN2(n1848), .Q(n4027) );
  NOR2X0 U5362 ( .IN1(n1585), .IN2(n4124), .QN(g23357) );
  XOR2X1 U5363 ( .IN1(n2484), .IN2(n4479), .Q(n4124) );
  INVX0 U5364 ( .IN(n2393), .QN(n2151) );
  INVX0 U5365 ( .IN(n2321), .QN(n2049) );
  INVX0 U5366 ( .IN(n2249), .QN(n1947) );
  INVX0 U5367 ( .IN(n2460), .QN(n1846) );
  INVX0 U5368 ( .IN(n2371), .QN(n2153) );
  INVX0 U5369 ( .IN(n2299), .QN(n2051) );
  INVX0 U5370 ( .IN(n2227), .QN(n1949) );
  INVX0 U5371 ( .IN(n2467), .QN(n1848) );
  INVX0 U5372 ( .IN(n3625), .QN(n2103) );
  INVX0 U5373 ( .IN(n3652), .QN(n2001) );
  INVX0 U5374 ( .IN(n3670), .QN(n1899) );
  INVX0 U5375 ( .IN(n3677), .QN(n1795) );
  INVX0 U5376 ( .IN(n3004), .QN(n2106) );
  INVX0 U5377 ( .IN(n3012), .QN(n2004) );
  INVX0 U5378 ( .IN(n3020), .QN(n1902) );
  INVX0 U5379 ( .IN(n3027), .QN(n1798) );
  NAND2X0 U5380 ( .IN1(n3713), .IN2(n3714), .QN(n3443) );
  NAND3X0 U5381 ( .IN1(n3449), .IN2(n3447), .IN3(n2110), .QN(n3713) );
  NAND3X0 U5382 ( .IN1(n1691), .IN2(n3448), .IN3(n2091), .QN(n3714) );
  NAND2X0 U5383 ( .IN1(n3719), .IN2(n3720), .QN(n3455) );
  NAND3X0 U5384 ( .IN1(n3461), .IN2(n3459), .IN3(n2007), .QN(n3719) );
  NAND3X0 U5385 ( .IN1(n1634), .IN2(n3460), .IN3(n1989), .QN(n3720) );
  NAND2X0 U5386 ( .IN1(n3725), .IN2(n3726), .QN(n3467) );
  NAND3X0 U5387 ( .IN1(n3473), .IN2(n3471), .IN3(n1905), .QN(n3725) );
  NAND3X0 U5388 ( .IN1(n1653), .IN2(n3472), .IN3(n1887), .QN(n3726) );
  NAND2X0 U5389 ( .IN1(n3730), .IN2(n3731), .QN(n3476) );
  NAND3X0 U5390 ( .IN1(n3482), .IN2(n3480), .IN3(n1801), .QN(n3730) );
  NAND3X0 U5391 ( .IN1(n1672), .IN2(n3481), .IN3(n1783), .QN(n3731) );
  INVX0 U5392 ( .IN(n3270), .QN(n2120) );
  INVX0 U5393 ( .IN(n3311), .QN(n2018) );
  INVX0 U5394 ( .IN(n3351), .QN(n1916) );
  INVX0 U5395 ( .IN(n3390), .QN(n1812) );
  INVX0 U5396 ( .IN(n2390), .QN(n2157) );
  INVX0 U5397 ( .IN(n2318), .QN(n2055) );
  INVX0 U5398 ( .IN(n2246), .QN(n1953) );
  INVX0 U5399 ( .IN(n2456), .QN(n1852) );
  INVX0 U5400 ( .IN(n2357), .QN(n2158) );
  INVX0 U5401 ( .IN(n2285), .QN(n2056) );
  INVX0 U5402 ( .IN(n2213), .QN(n1954) );
  INVX0 U5403 ( .IN(n2436), .QN(n1853) );
  INVX0 U5404 ( .IN(n3447), .QN(n2091) );
  INVX0 U5405 ( .IN(n3459), .QN(n1989) );
  INVX0 U5406 ( .IN(n3471), .QN(n1887) );
  INVX0 U5407 ( .IN(n3480), .QN(n1783) );
  INVX0 U5408 ( .IN(n2481), .QN(n1585) );
  INVX0 U5409 ( .IN(n3256), .QN(n1766) );
  INVX0 U5410 ( .IN(n3297), .QN(n1764) );
  INVX0 U5411 ( .IN(n3338), .QN(n1762) );
  INVX0 U5412 ( .IN(n3378), .QN(n1760) );
  XOR2X1 U5413 ( .IN1(n2998), .IN2(n4285), .Q(n2996) );
  NAND2X0 U5414 ( .IN1(n2999), .IN2(n3000), .QN(n2998) );
  OR4X1 U5415 ( .IN1(n2791), .IN2(n1693), .IN3(n2089), .IN4(n4285), .Q(n3000)
         );
  AO221X1 U5416 ( .IN1(n3001), .IN2(n2109), .IN3(n4285), .IN4(n3002), .IN5(
        n3003), .Q(n2999) );
  XOR2X1 U5417 ( .IN1(n3006), .IN2(n4284), .Q(n2997) );
  NAND2X0 U5418 ( .IN1(n3007), .IN2(n3008), .QN(n3006) );
  OR4X1 U5419 ( .IN1(n2610), .IN2(n1636), .IN3(n1987), .IN4(n4284), .Q(n3008)
         );
  AO221X1 U5420 ( .IN1(n3009), .IN2(n2008), .IN3(n4284), .IN4(n3010), .IN5(
        n3011), .Q(n3007) );
  XOR2X1 U5421 ( .IN1(n3021), .IN2(n4282), .Q(n3013) );
  NAND2X0 U5422 ( .IN1(n3022), .IN2(n3023), .QN(n3021) );
  OR4X1 U5423 ( .IN1(n2651), .IN2(n1674), .IN3(n1781), .IN4(n4282), .Q(n3023)
         );
  AO221X1 U5424 ( .IN1(n3024), .IN2(n1802), .IN3(n4282), .IN4(n3025), .IN5(
        n3026), .Q(n3022) );
  INVX0 U5425 ( .IN(n3257), .QN(n1765) );
  INVX0 U5426 ( .IN(n3298), .QN(n1763) );
  INVX0 U5427 ( .IN(n3339), .QN(n1761) );
  INVX0 U5428 ( .IN(n3379), .QN(n1759) );
  INVX0 U5429 ( .IN(n3702), .QN(n1748) );
  INVX0 U5430 ( .IN(n4201), .QN(n1629) );
  INVX0 U5431 ( .IN(n4212), .QN(n1628) );
  INVX0 U5432 ( .IN(n3003), .QN(n2090) );
  INVX0 U5433 ( .IN(n3011), .QN(n1988) );
  INVX0 U5434 ( .IN(n3019), .QN(n1886) );
  INVX0 U5435 ( .IN(n3026), .QN(n1782) );
  INVX0 U5436 ( .IN(n3174), .QN(n1829) );
  INVX0 U5437 ( .IN(n3706), .QN(n1747) );
  INVX0 U5438 ( .IN(n3700), .QN(n1574) );
  INVX0 U5439 ( .IN(n3935), .QN(n1626) );
  INVX0 U5440 ( .IN(n3449), .QN(n1691) );
  INVX0 U5441 ( .IN(n3461), .QN(n1634) );
  INVX0 U5442 ( .IN(n3473), .QN(n1653) );
  INVX0 U5443 ( .IN(n3482), .QN(n1672) );
  INVX0 U5444 ( .IN(n4659), .QN(n2126) );
  INVX0 U5445 ( .IN(n4657), .QN(n2024) );
  INVX0 U5446 ( .IN(n4655), .QN(n1922) );
  INVX0 U5447 ( .IN(n4653), .QN(n1820) );
  INVX0 U5448 ( .IN(n4660), .QN(n2125) );
  INVX0 U5449 ( .IN(n4658), .QN(n2023) );
  INVX0 U5450 ( .IN(n4656), .QN(n1921) );
  INVX0 U5451 ( .IN(n4654), .QN(n1819) );
  INVX0 U5452 ( .IN(n3951), .QN(n2146) );
  INVX0 U5453 ( .IN(n3954), .QN(n2145) );
  INVX0 U5454 ( .IN(n3971), .QN(n2044) );
  INVX0 U5455 ( .IN(n3974), .QN(n2043) );
  INVX0 U5456 ( .IN(n3991), .QN(n1942) );
  INVX0 U5457 ( .IN(n3996), .QN(n1941) );
  INVX0 U5458 ( .IN(n4013), .QN(n1841) );
  INVX0 U5459 ( .IN(n4014), .QN(n1840) );
  NOR2X0 U5460 ( .IN1(n4058), .IN2(n4305), .QN(n3736) );
  NOR2X0 U5461 ( .IN1(n4431), .IN2(n4123), .QN(n4059) );
  INVX0 U5462 ( .IN(n3950), .QN(n2147) );
  INVX0 U5463 ( .IN(n3953), .QN(n2045) );
  INVX0 U5464 ( .IN(n3973), .QN(n1943) );
  INVX0 U5465 ( .IN(n3993), .QN(n1842) );
  NOR2X0 U5466 ( .IN1(n4330), .IN2(n4423), .QN(n2486) );
  NOR2X0 U5467 ( .IN1(n4586), .IN2(n4423), .QN(g16802) );
  NOR2X0 U5468 ( .IN1(n3860), .IN2(n3734), .QN(g26037) );
  XOR2X1 U5469 ( .IN1(n3736), .IN2(n4291), .Q(n3860) );
  INVX0 U5470 ( .IN(n3678), .QN(n2164) );
  INVX0 U5471 ( .IN(n3486), .QN(n2062) );
  INVX0 U5472 ( .IN(n3490), .QN(n1960) );
  INVX0 U5473 ( .IN(n3494), .QN(n1859) );
  INVX0 U5474 ( .IN(n4170), .QN(n2086) );
  INVX0 U5475 ( .IN(n4172), .QN(n2084) );
  INVX0 U5476 ( .IN(n4173), .QN(n1984) );
  INVX0 U5477 ( .IN(n4175), .QN(n1982) );
  INVX0 U5478 ( .IN(n4176), .QN(n1882) );
  INVX0 U5479 ( .IN(n4178), .QN(n1880) );
  INVX0 U5480 ( .IN(n4179), .QN(n1778) );
  INVX0 U5481 ( .IN(n4180), .QN(n1776) );
  INVX0 U5482 ( .IN(n4362), .QN(n4690) );
  NAND2X0 U5483 ( .IN1(n1586), .IN2(n2485), .QN(n4274) );
  AO21X1 U5484 ( .IN1(n4423), .IN2(n4330), .IN3(n2486), .Q(n2485) );
  INVX0 U5485 ( .IN(n4153), .QN(n2162) );
  INVX0 U5486 ( .IN(n4159), .QN(n2060) );
  INVX0 U5487 ( .IN(n4165), .QN(n1958) );
  INVX0 U5488 ( .IN(n4168), .QN(n1857) );
  INVX0 U5489 ( .IN(n4200), .QN(n1579) );
  INVX0 U5490 ( .IN(n4147), .QN(n2148) );
  INVX0 U5491 ( .IN(n4151), .QN(n2046) );
  INVX0 U5492 ( .IN(n4157), .QN(n1944) );
  INVX0 U5493 ( .IN(n4163), .QN(n1843) );
  INVX0 U5494 ( .IN(n3855), .QN(n1828) );
  INVX0 U5495 ( .IN(n4146), .QN(n2165) );
  INVX0 U5496 ( .IN(n4150), .QN(n2063) );
  INVX0 U5497 ( .IN(n4156), .QN(n1961) );
  INVX0 U5498 ( .IN(n4162), .QN(n1860) );
  NOR2X0 U5499 ( .IN1(g499), .IN2(n4298), .QN(n2480) );
  NAND2X0 U5500 ( .IN1(n2478), .IN2(g499), .QN(n2439) );
  AO22X1 U5501 ( .IN1(g544), .IN2(g499), .IN3(n4206), .IN4(g548), .Q(g21851)
         );
  NOR2X0 U5502 ( .IN1(n4638), .IN2(g499), .QN(n4206) );
  NAND2X0 U5503 ( .IN1(n2426), .IN2(n2468), .QN(n4272) );
  AO221X1 U5504 ( .IN1(n1583), .IN2(DFF_449_n1), .IN3(n1832), .IN4(n2414), 
        .IN5(n1833), .Q(n2468) );
  AO221X1 U5505 ( .IN1(n1583), .IN2(DFF_448_n1), .IN3(n1832), .IN4(n2411), 
        .IN5(n1833), .Q(n2427) );
  AO222X1 U5506 ( .IN1(test_so22), .IN2(n2401), .IN3(n2402), .IN4(n1583), 
        .IN5(g557), .IN6(n2403), .Q(n4259) );
  NOR2X0 U5507 ( .IN1(n1833), .IN2(n2406), .QN(n2402) );
  XOR2X1 U5508 ( .IN1(n2404), .IN2(n2405), .Q(n2403) );
  XOR2X1 U5509 ( .IN1(n2407), .IN2(n2408), .Q(n2401) );
  NAND3X0 U5510 ( .IN1(n2434), .IN2(n2426), .IN3(n2435), .QN(n4266) );
  AO221X1 U5511 ( .IN1(n1583), .IN2(DFF_447_n1), .IN3(n1832), .IN4(n2409), 
        .IN5(n1833), .Q(n2435) );
  NAND3X0 U5512 ( .IN1(n2434), .IN2(n2426), .IN3(n2447), .QN(n4269) );
  AO221X1 U5513 ( .IN1(n1583), .IN2(DFF_444_n1), .IN3(n1832), .IN4(n2418), 
        .IN5(n1833), .Q(n2447) );
  NAND3X0 U5514 ( .IN1(n2440), .IN2(n2426), .IN3(n2441), .QN(n4267) );
  AO221X1 U5515 ( .IN1(n1583), .IN2(DFF_446_n1), .IN3(n1832), .IN4(n2413), 
        .IN5(n1833), .Q(n2441) );
  NAND3X0 U5516 ( .IN1(n2440), .IN2(n2426), .IN3(n2443), .QN(n4268) );
  AO221X1 U5517 ( .IN1(n1583), .IN2(DFF_445_n1), .IN3(n1832), .IN4(n2412), 
        .IN5(n1833), .Q(n2443) );
  AO21X1 U5518 ( .IN1(n2446), .IN2(n2405), .IN3(n2452), .Q(n4270) );
  OA221X1 U5519 ( .IN1(n2417), .IN2(n2453), .IN3(g537), .IN4(n2454), .IN5(
        n2455), .Q(n2452) );
  AO21X1 U5520 ( .IN1(n2446), .IN2(n2404), .IN3(n2461), .Q(n4271) );
  OA221X1 U5521 ( .IN1(n2416), .IN2(n2453), .IN3(g536), .IN4(n2454), .IN5(
        n2455), .Q(n2461) );
  AO21X1 U5522 ( .IN1(g2631), .IN2(n4303), .IN3(n2400), .Q(n2363) );
  AO21X1 U5523 ( .IN1(g1937), .IN2(n4297), .IN3(n2328), .Q(n2291) );
  AO21X1 U5524 ( .IN1(g1243), .IN2(n4304), .IN3(n2256), .Q(n2219) );
  AO21X1 U5525 ( .IN1(g557), .IN2(n4310), .IN3(n2479), .Q(n2453) );
  AO21X1 U5526 ( .IN1(g2584), .IN2(n4352), .IN3(n2400), .Q(n2365) );
  AO21X1 U5527 ( .IN1(g1890), .IN2(n4311), .IN3(n2328), .Q(n2293) );
  AO21X1 U5528 ( .IN1(g1196), .IN2(n4353), .IN3(n2256), .Q(n2221) );
  AO21X1 U5529 ( .IN1(test_so22), .IN2(n4360), .IN3(n2479), .Q(n2455) );
  NAND2X0 U5530 ( .IN1(n2347), .IN2(n2378), .QN(n4256) );
  AO221X1 U5531 ( .IN1(n1570), .IN2(DFF_1499_n1), .IN3(n2136), .IN4(n2342), 
        .IN5(n2137), .Q(n2378) );
  NAND2X0 U5532 ( .IN1(n2347), .IN2(n2348), .QN(n4251) );
  AO221X1 U5533 ( .IN1(n1570), .IN2(DFF_1498_n1), .IN3(n2136), .IN4(n2339), 
        .IN5(n2137), .Q(n2348) );
  NAND2X0 U5534 ( .IN1(n2275), .IN2(n2306), .QN(n4247) );
  AO221X1 U5535 ( .IN1(n1568), .IN2(DFF_1149_n1), .IN3(n2034), .IN4(n2270), 
        .IN5(n2035), .Q(n2306) );
  NAND2X0 U5536 ( .IN1(n2275), .IN2(n2276), .QN(n4242) );
  AO221X1 U5537 ( .IN1(n1568), .IN2(DFF_1148_n1), .IN3(n2034), .IN4(n2267), 
        .IN5(n2035), .Q(n2276) );
  NAND2X0 U5538 ( .IN1(n2203), .IN2(n2234), .QN(n4238) );
  AO221X1 U5539 ( .IN1(n1566), .IN2(DFF_799_n1), .IN3(n1932), .IN4(n2198), 
        .IN5(n1933), .Q(n2234) );
  NAND2X0 U5540 ( .IN1(n2203), .IN2(n2204), .QN(n4233) );
  AO221X1 U5541 ( .IN1(n1566), .IN2(DFF_798_n1), .IN3(n1932), .IN4(n2195), 
        .IN5(n1933), .Q(n2204) );
  AND3X1 U5542 ( .IN1(n4303), .IN2(n4352), .IN3(g2599), .Q(n2400) );
  AND3X1 U5543 ( .IN1(n4297), .IN2(n4311), .IN3(g1905), .Q(n2328) );
  AND3X1 U5544 ( .IN1(n4304), .IN2(n4353), .IN3(g1211), .Q(n2256) );
  AND3X1 U5545 ( .IN1(n4310), .IN2(n4360), .IN3(g525), .Q(n2479) );
  NAND3X0 U5546 ( .IN1(n2355), .IN2(n2347), .IN3(n2356), .QN(n4252) );
  AO221X1 U5547 ( .IN1(n1570), .IN2(DFF_1497_n1), .IN3(n2136), .IN4(n2337), 
        .IN5(n2137), .Q(n2356) );
  NAND3X0 U5548 ( .IN1(n2355), .IN2(n2347), .IN3(n2372), .QN(n4254) );
  AO221X1 U5549 ( .IN1(n1570), .IN2(DFF_1494_n1), .IN3(n2136), .IN4(n2340), 
        .IN5(n2137), .Q(n2372) );
  NAND3X0 U5550 ( .IN1(n2283), .IN2(n2275), .IN3(n2284), .QN(n4243) );
  AO221X1 U5551 ( .IN1(n1568), .IN2(DFF_1147_n1), .IN3(n2034), .IN4(n2265), 
        .IN5(n2035), .Q(n2284) );
  NAND3X0 U5552 ( .IN1(n2283), .IN2(n2275), .IN3(n2300), .QN(n4245) );
  AO221X1 U5553 ( .IN1(n1568), .IN2(DFF_1144_n1), .IN3(n2034), .IN4(n2268), 
        .IN5(n2035), .Q(n2300) );
  NAND3X0 U5554 ( .IN1(n2211), .IN2(n2203), .IN3(n2212), .QN(n4234) );
  AO221X1 U5555 ( .IN1(n1566), .IN2(DFF_797_n1), .IN3(n1932), .IN4(n2193), 
        .IN5(n1933), .Q(n2212) );
  NAND3X0 U5556 ( .IN1(n2211), .IN2(n2203), .IN3(n2228), .QN(n4236) );
  AO221X1 U5557 ( .IN1(n1566), .IN2(DFF_794_n1), .IN3(n1932), .IN4(n2196), 
        .IN5(n1933), .Q(n2228) );
  NAND3X0 U5558 ( .IN1(n2375), .IN2(n2347), .IN3(n2376), .QN(n4255) );
  AO221X1 U5559 ( .IN1(n1570), .IN2(DFF_1496_n1), .IN3(n2136), .IN4(n2344), 
        .IN5(n2137), .Q(n2376) );
  NAND3X0 U5560 ( .IN1(n2375), .IN2(n2347), .IN3(n2383), .QN(n4257) );
  AO221X1 U5561 ( .IN1(n1570), .IN2(DFF_1495_n1), .IN3(n2136), .IN4(n2346), 
        .IN5(n2137), .Q(n2383) );
  NAND3X0 U5562 ( .IN1(n2303), .IN2(n2275), .IN3(n2304), .QN(n4246) );
  AO221X1 U5563 ( .IN1(n1568), .IN2(DFF_1146_n1), .IN3(n2034), .IN4(n2272), 
        .IN5(n2035), .Q(n2304) );
  NAND3X0 U5564 ( .IN1(n2303), .IN2(n2275), .IN3(n2311), .QN(n4248) );
  AO221X1 U5565 ( .IN1(n1568), .IN2(DFF_1145_n1), .IN3(n2034), .IN4(n2274), 
        .IN5(n2035), .Q(n2311) );
  NAND3X0 U5566 ( .IN1(n2231), .IN2(n2203), .IN3(n2232), .QN(n4237) );
  AO221X1 U5567 ( .IN1(n1566), .IN2(DFF_796_n1), .IN3(n1932), .IN4(n2200), 
        .IN5(n1933), .Q(n2232) );
  NAND3X0 U5568 ( .IN1(n2231), .IN2(n2203), .IN3(n2239), .QN(n4239) );
  AO221X1 U5569 ( .IN1(n1566), .IN2(DFF_795_n1), .IN3(n1932), .IN4(n2202), 
        .IN5(n1933), .Q(n2239) );
  NOR3X0 U5570 ( .IN1(g2637), .IN2(g2633), .IN3(g30072), .QN(n2385) );
  NOR3X0 U5571 ( .IN1(g1249), .IN2(g1245), .IN3(n1817), .QN(n2241) );
  NAND2X0 U5572 ( .IN1(n2385), .IN2(g2574), .QN(n2360) );
  NAND2X0 U5573 ( .IN1(n2241), .IN2(g1186), .QN(n2216) );
  NOR4X0 U5574 ( .IN1(g3013), .IN2(g3024), .IN3(test_so98), .IN4(n4221), .QN(
        n4144) );
  OR2X1 U5575 ( .IN1(g3006), .IN2(g3002), .Q(n4221) );
  OA222X1 U5576 ( .IN1(n4524), .IN2(g2391), .IN3(n4509), .IN4(g2392), .IN5(
        n4516), .IN6(g2390), .Q(n2778) );
  OA222X1 U5577 ( .IN1(n4525), .IN2(g1697), .IN3(n4511), .IN4(g1698), .IN5(
        n4518), .IN6(g1696), .Q(n2597) );
  OA222X1 U5578 ( .IN1(n4676), .IN2(test_so18), .IN3(n4506), .IN4(g317), .IN5(
        n4520), .IN6(g315), .Q(n2638) );
  AO21X1 U5579 ( .IN1(n2361), .IN2(n2332), .IN3(n2389), .Q(n4258) );
  OA221X1 U5580 ( .IN1(n2345), .IN2(n2363), .IN3(g2611), .IN4(n2364), .IN5(
        n2365), .Q(n2389) );
  AO21X1 U5581 ( .IN1(n2361), .IN2(n2333), .IN3(n2362), .Q(n4253) );
  OA221X1 U5582 ( .IN1(n2341), .IN2(n2363), .IN3(test_so91), .IN4(n2364), 
        .IN5(n2365), .Q(n2362) );
  AO21X1 U5583 ( .IN1(n2289), .IN2(n2260), .IN3(n2317), .Q(n4249) );
  OA221X1 U5584 ( .IN1(n2273), .IN2(n2291), .IN3(g1917), .IN4(n2292), .IN5(
        n2293), .Q(n2317) );
  AO21X1 U5585 ( .IN1(n2289), .IN2(n2261), .IN3(n2290), .Q(n4244) );
  OA221X1 U5586 ( .IN1(n2269), .IN2(n2291), .IN3(g1916), .IN4(n2292), .IN5(
        n2293), .Q(n2290) );
  AO21X1 U5587 ( .IN1(n2217), .IN2(n2188), .IN3(n2245), .Q(n4240) );
  OA221X1 U5588 ( .IN1(n2201), .IN2(n2219), .IN3(g1223), .IN4(n2220), .IN5(
        n2221), .Q(n2245) );
  AO21X1 U5589 ( .IN1(n2217), .IN2(n2189), .IN3(n2218), .Q(n4235) );
  OA221X1 U5590 ( .IN1(n2197), .IN2(n2219), .IN3(g1222), .IN4(n2220), .IN5(
        n2221), .Q(n2218) );
  OA222X1 U5591 ( .IN1(n4524), .IN2(g2388), .IN3(n4509), .IN4(g2389), .IN5(
        n4516), .IN6(g2387), .Q(n4116) );
  OA222X1 U5592 ( .IN1(n4525), .IN2(g1694), .IN3(n4511), .IN4(g1695), .IN5(
        n4518), .IN6(g1693), .Q(n4117) );
  OA222X1 U5593 ( .IN1(n4676), .IN2(g313), .IN3(n4506), .IN4(g314), .IN5(n4520), .IN6(g312), .Q(n4119) );
  OA222X1 U5594 ( .IN1(n4359), .IN2(g724), .IN3(n4295), .IN4(g722), .IN5(n4309), .IN6(g723), .Q(n2460) );
  OA222X1 U5595 ( .IN1(n4356), .IN2(g2798), .IN3(n4292), .IN4(test_so94), 
        .IN5(n4306), .IN6(g2797), .Q(n2393) );
  OA222X1 U5596 ( .IN1(n4357), .IN2(g2104), .IN3(n4293), .IN4(g2102), .IN5(
        n4307), .IN6(g2103), .Q(n2321) );
  OA222X1 U5597 ( .IN1(n4358), .IN2(g1410), .IN3(n4294), .IN4(g1408), .IN5(
        n4308), .IN6(g1409), .Q(n2249) );
  OA222X1 U5598 ( .IN1(n4359), .IN2(test_so30), .IN3(n4295), .IN4(g725), .IN5(
        n4309), .IN6(g726), .Q(n2467) );
  OA222X1 U5599 ( .IN1(n4356), .IN2(g2801), .IN3(n4292), .IN4(g2799), .IN5(
        n4306), .IN6(g2800), .Q(n2371) );
  OA222X1 U5600 ( .IN1(n4357), .IN2(test_so72), .IN3(n4293), .IN4(g2105), 
        .IN5(n4307), .IN6(g2106), .Q(n2299) );
  OA222X1 U5601 ( .IN1(n4358), .IN2(g1413), .IN3(n4294), .IN4(g1411), .IN5(
        n4308), .IN6(g1412), .Q(n2227) );
  AO222X1 U5602 ( .IN1(g2300), .IN2(g7084), .IN3(g2303), .IN4(n4679), .IN5(
        g2297), .IN6(g2214), .Q(n2500) );
  AO222X1 U5603 ( .IN1(g2309), .IN2(g7084), .IN3(g2312), .IN4(n4679), .IN5(
        g2306), .IN6(g2214), .Q(n2512) );
  AO222X1 U5604 ( .IN1(test_so56), .IN2(n4589), .IN3(g1609), .IN4(n4684), 
        .IN5(g1603), .IN6(g1520), .Q(n2527) );
  AO222X1 U5605 ( .IN1(g1615), .IN2(g6782), .IN3(g1618), .IN4(n4684), .IN5(
        g1612), .IN6(g1520), .Q(n2538) );
  AO222X1 U5606 ( .IN1(g225), .IN2(g6313), .IN3(g228), .IN4(n4694), .IN5(g222), 
        .IN6(g138), .Q(n2579) );
  AO222X1 U5607 ( .IN1(g234), .IN2(g6313), .IN3(g237), .IN4(n4694), .IN5(g231), 
        .IN6(g138), .Q(n2590) );
  OA222X1 U5608 ( .IN1(n4356), .IN2(g2777), .IN3(n4292), .IN4(g2775), .IN5(
        n4306), .IN6(g2776), .Q(n2368) );
  OA222X1 U5609 ( .IN1(n4357), .IN2(g2083), .IN3(n4293), .IN4(g2081), .IN5(
        n4307), .IN6(g2082), .Q(n2296) );
  OA222X1 U5610 ( .IN1(n4358), .IN2(g1389), .IN3(n4294), .IN4(g1387), .IN5(
        n4308), .IN6(g1388), .Q(n2224) );
  OA222X1 U5611 ( .IN1(n4356), .IN2(g2783), .IN3(n4292), .IN4(test_so93), 
        .IN5(n4306), .IN6(g2782), .Q(n2352) );
  OA222X1 U5612 ( .IN1(n4356), .IN2(g2780), .IN3(n4292), .IN4(g2778), .IN5(
        n4306), .IN6(g2779), .Q(n2382) );
  OA222X1 U5613 ( .IN1(n4357), .IN2(g2089), .IN3(n4293), .IN4(g2087), .IN5(
        n4307), .IN6(g2088), .Q(n2280) );
  OA222X1 U5614 ( .IN1(n4357), .IN2(g2086), .IN3(n4293), .IN4(g2084), .IN5(
        n4307), .IN6(g2085), .Q(n2310) );
  OA222X1 U5615 ( .IN1(n4358), .IN2(g1395), .IN3(n4294), .IN4(g1393), .IN5(
        n4308), .IN6(g1394), .Q(n2208) );
  OA222X1 U5616 ( .IN1(n4358), .IN2(g1392), .IN3(n4294), .IN4(g1390), .IN5(
        n4308), .IN6(g1391), .Q(n2238) );
  OA222X1 U5617 ( .IN1(n4359), .IN2(g706), .IN3(n4295), .IN4(g704), .IN5(n4309), .IN6(g705), .Q(n2471) );
  OA222X1 U5618 ( .IN1(n4359), .IN2(g703), .IN3(n4295), .IN4(g701), .IN5(n4309), .IN6(g702), .Q(n2464) );
  OA222X1 U5619 ( .IN1(n4359), .IN2(g709), .IN3(n4295), .IN4(g707), .IN5(n4309), .IN6(g708), .Q(n2431) );
  OA222X1 U5620 ( .IN1(n4359), .IN2(g700), .IN3(n4295), .IN4(g698), .IN5(n4309), .IN6(g699), .Q(n2456) );
  OA222X1 U5621 ( .IN1(n4356), .IN2(g2774), .IN3(n4292), .IN4(g2772), .IN5(
        n4306), .IN6(g2773), .Q(n2390) );
  OA222X1 U5622 ( .IN1(n4357), .IN2(g2080), .IN3(n4293), .IN4(g2078), .IN5(
        n4307), .IN6(g2079), .Q(n2318) );
  OA222X1 U5623 ( .IN1(n4358), .IN2(g1386), .IN3(n4294), .IN4(g1384), .IN5(
        n4308), .IN6(test_so49), .Q(n2246) );
  OA222X1 U5624 ( .IN1(n4359), .IN2(g712), .IN3(n4295), .IN4(g710), .IN5(n4309), .IN6(test_so29), .Q(n2436) );
  OA222X1 U5625 ( .IN1(n4356), .IN2(g2786), .IN3(n4292), .IN4(g2784), .IN5(
        n4306), .IN6(g2785), .Q(n2357) );
  OA222X1 U5626 ( .IN1(n4357), .IN2(test_so71), .IN3(n4293), .IN4(g2090), 
        .IN5(n4307), .IN6(g2091), .Q(n2285) );
  OA222X1 U5627 ( .IN1(n4358), .IN2(g1398), .IN3(n4294), .IN4(g1396), .IN5(
        n4308), .IN6(g1397), .Q(n2213) );
  AO222X1 U5628 ( .IN1(g2273), .IN2(n4587), .IN3(g2276), .IN4(n4679), .IN5(
        g2270), .IN6(g6837), .Q(n2498) );
  AO222X1 U5629 ( .IN1(g1579), .IN2(g6782), .IN3(g1582), .IN4(n4684), .IN5(
        g1576), .IN6(g6573), .Q(n2525) );
  AO222X1 U5630 ( .IN1(g198), .IN2(n4593), .IN3(g201), .IN4(n4694), .IN5(g195), 
        .IN6(g6231), .Q(n2577) );
  AND3X1 U5631 ( .IN1(n2982), .IN2(n3157), .IN3(n3158), .Q(g29112) );
  AND3X1 U5632 ( .IN1(n2985), .IN2(n3161), .IN3(n3162), .Q(g29111) );
  AND3X1 U5633 ( .IN1(n2988), .IN2(n3165), .IN3(n3166), .Q(g29110) );
  AND3X1 U5634 ( .IN1(n2991), .IN2(n3169), .IN3(n3170), .Q(g29109) );
  OA222X1 U5635 ( .IN1(n4356), .IN2(g2795), .IN3(n4292), .IN4(g2793), .IN5(
        n4306), .IN6(g2794), .Q(n2373) );
  OA222X1 U5636 ( .IN1(n4356), .IN2(g2792), .IN3(n4292), .IN4(g2790), .IN5(
        n4306), .IN6(g2791), .Q(n2384) );
  OA222X1 U5637 ( .IN1(n4357), .IN2(g2101), .IN3(n4293), .IN4(g2099), .IN5(
        n4307), .IN6(g2100), .Q(n2301) );
  OA222X1 U5638 ( .IN1(n4357), .IN2(g2098), .IN3(n4293), .IN4(g2096), .IN5(
        n4307), .IN6(g2097), .Q(n2312) );
  OA222X1 U5639 ( .IN1(n4358), .IN2(g1407), .IN3(n4294), .IN4(g1405), .IN5(
        n4308), .IN6(g1406), .Q(n2229) );
  OA222X1 U5640 ( .IN1(n4358), .IN2(g1404), .IN3(n4294), .IN4(g1402), .IN5(
        n4308), .IN6(g1403), .Q(n2240) );
  OA222X1 U5641 ( .IN1(n4359), .IN2(g721), .IN3(n4295), .IN4(g719), .IN5(n4309), .IN6(g720), .Q(n2448) );
  OA222X1 U5642 ( .IN1(n4359), .IN2(g718), .IN3(n4295), .IN4(g716), .IN5(n4309), .IN6(g717), .Q(n2444) );
  OA222X1 U5643 ( .IN1(n4359), .IN2(g715), .IN3(n4295), .IN4(g713), .IN5(n4309), .IN6(g714), .Q(n2442) );
  OA222X1 U5644 ( .IN1(n4356), .IN2(g2789), .IN3(n4292), .IN4(g2787), .IN5(
        n4306), .IN6(g2788), .Q(n2377) );
  OA222X1 U5645 ( .IN1(n4357), .IN2(g2095), .IN3(n4293), .IN4(g2093), .IN5(
        n4307), .IN6(g2094), .Q(n2305) );
  OA222X1 U5646 ( .IN1(n4358), .IN2(test_so50), .IN3(n4294), .IN4(g1399), 
        .IN5(n4308), .IN6(g1400), .Q(n2233) );
  AO21X1 U5647 ( .IN1(n4121), .IN2(n1582), .IN3(n1581), .Q(n2422) );
  NAND4X0 U5648 ( .IN1(g3032), .IN2(g3018), .IN3(n4350), .IN4(n4480), .QN(
        n4121) );
  AND3X1 U5649 ( .IN1(n4064), .IN2(n3742), .IN3(n1581), .Q(g25191) );
  AO21X1 U5650 ( .IN1(g1880), .IN2(DFF_1099_n1), .IN3(n3155), .Q(n2961) );
  OA221X1 U5651 ( .IN1(g7052), .IN2(DFF_1100_n1), .IN3(n3156), .IN4(n4296), 
        .IN5(n4545), .Q(n3155) );
  AO222X1 U5652 ( .IN1(g2291), .IN2(n4587), .IN3(g2294), .IN4(n4679), .IN5(
        g2288), .IN6(g6837), .Q(n2501) );
  AO222X1 U5653 ( .IN1(g1597), .IN2(n4589), .IN3(g1600), .IN4(n4684), .IN5(
        g1594), .IN6(g6573), .Q(n2528) );
  AO222X1 U5654 ( .IN1(g216), .IN2(n4593), .IN3(g219), .IN4(n4694), .IN5(g213), 
        .IN6(g6231), .Q(n2580) );
  AO222X1 U5655 ( .IN1(g2336), .IN2(g7084), .IN3(g2339), .IN4(n4679), .IN5(
        g2333), .IN6(g2214), .Q(n2502) );
  AO222X1 U5656 ( .IN1(g1642), .IN2(n4589), .IN3(g1645), .IN4(n4684), .IN5(
        g1639), .IN6(g1520), .Q(n2529) );
  AO222X1 U5657 ( .IN1(g261), .IN2(g6313), .IN3(g264), .IN4(n4694), .IN5(g258), 
        .IN6(g138), .Q(n2581) );
  AOI222X1 U5658 ( .IN1(g2282), .IN2(g7084), .IN3(g2285), .IN4(n4679), .IN5(
        g2279), .IN6(g2214), .QN(n2511) );
  AOI222X1 U5659 ( .IN1(g1588), .IN2(g6782), .IN3(g1591), .IN4(n4684), .IN5(
        g1585), .IN6(g1520), .QN(n2537) );
  AOI222X1 U5660 ( .IN1(g207), .IN2(g6313), .IN3(g210), .IN4(n4694), .IN5(g204), .IN6(g138), .QN(n2589) );
  OA222X1 U5661 ( .IN1(n4359), .IN2(g733), .IN3(n4295), .IN4(g731), .IN5(n4309), .IN6(g732), .Q(n2475) );
  OA222X1 U5662 ( .IN1(n4356), .IN2(g2807), .IN3(n4292), .IN4(g2805), .IN5(
        n4306), .IN6(g2806), .Q(n2397) );
  OA222X1 U5663 ( .IN1(n4357), .IN2(g2113), .IN3(n4293), .IN4(g2111), .IN5(
        n4307), .IN6(g2112), .Q(n2325) );
  OA222X1 U5664 ( .IN1(n4358), .IN2(g1419), .IN3(n4294), .IN4(g1417), .IN5(
        n4308), .IN6(g1418), .Q(n2253) );
  NAND2X0 U5665 ( .IN1(n2425), .IN2(g3028), .QN(n4102) );
  AND3X1 U5666 ( .IN1(n4128), .IN2(n4066), .IN3(n1581), .Q(g23330) );
  AO222X1 U5667 ( .IN1(g1196), .IN2(n2185), .IN3(n2186), .IN4(n1566), .IN5(
        g1243), .IN6(n2187), .Q(n4232) );
  NOR2X0 U5668 ( .IN1(n1933), .IN2(n2190), .QN(n2186) );
  XOR2X1 U5669 ( .IN1(n2188), .IN2(n2189), .Q(n2187) );
  XOR2X1 U5670 ( .IN1(n2191), .IN2(n2192), .Q(n2185) );
  AND4X1 U5671 ( .IN1(g3028), .IN2(g3018), .IN3(n4207), .IN4(n4129), .Q(n4553)
         );
  OA221X1 U5672 ( .IN1(g7302), .IN2(DFF_1450_n1), .IN3(n2961), .IN4(n4314), 
        .IN5(n4543), .Q(n2960) );
  AO22X1 U5673 ( .IN1(g2733), .IN2(n4292), .IN3(n4144), .IN4(g2703), .Q(g20375) );
  AO22X1 U5674 ( .IN1(g2039), .IN2(n4293), .IN3(n4144), .IN4(g2009), .Q(g20353) );
  AO22X1 U5675 ( .IN1(g1345), .IN2(n4294), .IN3(n4144), .IN4(g1315), .Q(g20333) );
  AO22X1 U5676 ( .IN1(g659), .IN2(n4295), .IN3(n4144), .IN4(g629), .Q(g20314)
         );
  AO22X1 U5677 ( .IN1(g2628), .IN2(n4299), .IN3(n4600), .IN4(n4662), .Q(g21847) );
  AO22X1 U5678 ( .IN1(g1934), .IN2(n4366), .IN3(n4612), .IN4(n4661), .Q(g21845) );
  AO22X1 U5679 ( .IN1(g554), .IN2(n4313), .IN3(n4634), .IN4(n4661), .Q(g21842)
         );
  AO22X1 U5680 ( .IN1(g1240), .IN2(n4300), .IN3(n4624), .IN4(n4661), .Q(g21843) );
  AO22X1 U5681 ( .IN1(g2348), .IN2(n4680), .IN3(n2657), .IN4(g2241), .Q(g30694) );
  AO22X1 U5682 ( .IN1(g1654), .IN2(n4685), .IN3(n2664), .IN4(g1547), .Q(g30689) );
  AO22X1 U5683 ( .IN1(g273), .IN2(n4695), .IN3(n2693), .IN4(g165), .Q(g30675)
         );
  AO22X1 U5684 ( .IN1(g2342), .IN2(n4683), .IN3(n2657), .IN4(g2214), .Q(g30686) );
  AO22X1 U5685 ( .IN1(g2297), .IN2(n4683), .IN3(g6837), .IN4(n2711), .Q(g30652) );
  AO22X1 U5686 ( .IN1(g1648), .IN2(n4317), .IN3(n2664), .IN4(g1520), .Q(g30678) );
  AO22X1 U5687 ( .IN1(g1603), .IN2(n4317), .IN3(g6573), .IN4(n2730), .Q(g30644) );
  AO22X1 U5688 ( .IN1(g267), .IN2(n4318), .IN3(n2693), .IN4(g138), .Q(g30661)
         );
  AO22X1 U5689 ( .IN1(g222), .IN2(n4318), .IN3(g6231), .IN4(n2762), .Q(g30635)
         );
  AO22X1 U5690 ( .IN1(g2345), .IN2(n4682), .IN3(n2657), .IN4(g7084), .Q(g30691) );
  AO22X1 U5691 ( .IN1(g2300), .IN2(n4681), .IN3(n4587), .IN4(n2711), .Q(g30659) );
  AO22X1 U5692 ( .IN1(g1651), .IN2(n4686), .IN3(n2664), .IN4(n4589), .Q(g30684) );
  AO22X1 U5693 ( .IN1(test_so56), .IN2(n4686), .IN3(g6782), .IN4(n2730), .Q(
        g30650) );
  AO22X1 U5694 ( .IN1(g270), .IN2(n4696), .IN3(n2693), .IN4(g6313), .Q(g30669)
         );
  AO22X1 U5695 ( .IN1(g225), .IN2(n4696), .IN3(n4593), .IN4(n2762), .Q(g30636)
         );
  AO22X1 U5696 ( .IN1(g2661), .IN2(n4314), .IN3(n4075), .IN4(n4604), .Q(g24527) );
  AO22X1 U5697 ( .IN1(g1967), .IN2(n4296), .IN3(n4079), .IN4(n4616), .Q(g24513) );
  AO22X1 U5698 ( .IN1(g1273), .IN2(n4371), .IN3(n4085), .IN4(n4628), .Q(g24501) );
  AO22X1 U5699 ( .IN1(g587), .IN2(n4298), .IN3(n4091), .IN4(n4638), .Q(g24491)
         );
  AO22X1 U5700 ( .IN1(g2685), .IN2(n4299), .IN3(n4600), .IN4(n3249), .Q(g28367) );
  AO22X1 U5701 ( .IN1(g2694), .IN2(n4299), .IN3(n4600), .IN4(n3248), .Q(g28371) );
  AO22X1 U5702 ( .IN1(g2676), .IN2(n4299), .IN3(n4074), .IN4(n4600), .Q(g24557) );
  AO22X1 U5703 ( .IN1(g2667), .IN2(n4299), .IN3(n4075), .IN4(n4600), .Q(g24547) );
  AO22X1 U5704 ( .IN1(g1991), .IN2(n4366), .IN3(n4612), .IN4(n3258), .Q(g28361) );
  AO22X1 U5705 ( .IN1(g2000), .IN2(n4366), .IN3(n4612), .IN4(n3250), .Q(g28366) );
  AO22X1 U5706 ( .IN1(g1982), .IN2(n4366), .IN3(n4076), .IN4(n4612), .Q(g24545) );
  AO22X1 U5707 ( .IN1(g1973), .IN2(n4366), .IN3(n4079), .IN4(n4612), .Q(g24534) );
  AO22X1 U5708 ( .IN1(g1297), .IN2(n4300), .IN3(n4624), .IN4(n3299), .Q(g28354) );
  AO22X1 U5709 ( .IN1(g1306), .IN2(n4300), .IN3(n4624), .IN4(n3259), .Q(g28360) );
  AO22X1 U5710 ( .IN1(g1288), .IN2(n4300), .IN3(n4080), .IN4(n4624), .Q(g24532) );
  AO22X1 U5711 ( .IN1(g1279), .IN2(n4300), .IN3(n4085), .IN4(n4624), .Q(g24521) );
  AO22X1 U5712 ( .IN1(g611), .IN2(n4313), .IN3(n4634), .IN4(n3340), .Q(g28348)
         );
  AO22X1 U5713 ( .IN1(test_so26), .IN2(n4313), .IN3(n4634), .IN4(n3300), .Q(
        g28353) );
  AO22X1 U5714 ( .IN1(g602), .IN2(n4313), .IN3(n4086), .IN4(n4634), .Q(g24519)
         );
  AO22X1 U5715 ( .IN1(g593), .IN2(n4313), .IN3(n4091), .IN4(n4634), .Q(g24507)
         );
  AO22X1 U5716 ( .IN1(g2670), .IN2(n4314), .IN3(n4074), .IN4(g7302), .Q(g24538) );
  AO22X1 U5717 ( .IN1(g1976), .IN2(n4296), .IN3(n4076), .IN4(g7052), .Q(g24525) );
  AO22X1 U5718 ( .IN1(g1282), .IN2(n4371), .IN3(n4080), .IN4(g6750), .Q(g24511) );
  AO22X1 U5719 ( .IN1(g596), .IN2(n4298), .IN3(n4086), .IN4(g6485), .Q(g24499)
         );
  AO22X1 U5720 ( .IN1(g2303), .IN2(n4680), .IN3(g2241), .IN4(n2711), .Q(g30665) );
  AO22X1 U5721 ( .IN1(g1609), .IN2(n4685), .IN3(g1547), .IN4(n2730), .Q(g30656) );
  AO22X1 U5722 ( .IN1(g228), .IN2(n4695), .IN3(g165), .IN4(n2762), .Q(g30639)
         );
  AO22X1 U5723 ( .IN1(g605), .IN2(n4298), .IN3(g6485), .IN4(n3340), .Q(g28342)
         );
  AO22X1 U5724 ( .IN1(g614), .IN2(n4298), .IN3(n4638), .IN4(n3300), .Q(g28345)
         );
  AO22X1 U5725 ( .IN1(test_so90), .IN2(n4370), .IN3(n4602), .IN4(n3249), .Q(
        g28363) );
  AO22X1 U5726 ( .IN1(g2673), .IN2(n4370), .IN3(n4074), .IN4(n4602), .Q(g24548) );
  AO22X1 U5727 ( .IN1(g2664), .IN2(n4370), .IN3(n4075), .IN4(n4602), .Q(g24537) );
  AO22X1 U5728 ( .IN1(g2679), .IN2(n4314), .IN3(g7302), .IN4(n3249), .Q(g28358) );
  AO22X1 U5729 ( .IN1(g2691), .IN2(n4370), .IN3(n4602), .IN4(n3248), .Q(g28368) );
  AO22X1 U5730 ( .IN1(g2688), .IN2(n4314), .IN3(n4604), .IN4(n3248), .Q(g28364) );
  AO22X1 U5731 ( .IN1(g1988), .IN2(n4315), .IN3(n4614), .IN4(n3258), .Q(g28356) );
  AO22X1 U5732 ( .IN1(g1970), .IN2(n4315), .IN3(n4079), .IN4(n4614), .Q(g24524) );
  AO22X1 U5733 ( .IN1(g1985), .IN2(n4296), .IN3(g7052), .IN4(n3258), .Q(g28352) );
  AO22X1 U5734 ( .IN1(g1997), .IN2(n4315), .IN3(n4614), .IN4(n3250), .Q(g28362) );
  AO22X1 U5735 ( .IN1(g1979), .IN2(n4315), .IN3(n4076), .IN4(n4614), .Q(g24535) );
  AO22X1 U5736 ( .IN1(g1994), .IN2(n4296), .IN3(n4616), .IN4(n3250), .Q(g28357) );
  AO22X1 U5737 ( .IN1(g1294), .IN2(n4316), .IN3(n4626), .IN4(n3299), .Q(g28350) );
  AO22X1 U5738 ( .IN1(g1291), .IN2(n4371), .IN3(g6750), .IN4(n3299), .Q(g28346) );
  AO22X1 U5739 ( .IN1(g1303), .IN2(n4316), .IN3(n4626), .IN4(n3259), .Q(g28355) );
  AO22X1 U5740 ( .IN1(g1285), .IN2(n4316), .IN3(n4080), .IN4(n4626), .Q(g24522) );
  AO22X1 U5741 ( .IN1(g1276), .IN2(n4316), .IN3(n4085), .IN4(n4626), .Q(g24510) );
  AO22X1 U5742 ( .IN1(g1300), .IN2(n4371), .IN3(n4628), .IN4(n3259), .Q(g28351) );
  AO22X1 U5743 ( .IN1(g599), .IN2(n4372), .IN3(n4086), .IN4(n4636), .Q(g24508)
         );
  AO22X1 U5744 ( .IN1(g590), .IN2(n4372), .IN3(n4091), .IN4(n4636), .Q(g24498)
         );
  AO22X1 U5745 ( .IN1(g608), .IN2(n4372), .IN3(n4636), .IN4(n3340), .Q(g28344)
         );
  AO22X1 U5746 ( .IN1(g617), .IN2(n4372), .IN3(n4636), .IN4(n3300), .Q(g28349)
         );
  AND4X1 U5747 ( .IN1(g3013), .IN2(g3002), .IN3(g3024), .IN4(n4208), .Q(n4129)
         );
  NOR4X0 U5748 ( .IN1(test_so98), .IN2(g3006), .IN3(g2993), .IN4(n4354), .QN(
        n4208) );
  ISOLANDX1 U5749 ( .D(g2133), .ISO(n3160), .Q(n3159) );
  ISOLANDX1 U5750 ( .D(g1439), .ISO(n3164), .Q(n3163) );
  ISOLANDX1 U5751 ( .D(g753), .ISO(n3168), .Q(n3167) );
  ISOLANDX1 U5752 ( .D(g65), .ISO(n3172), .Q(n3171) );
  ISOLANDX1 U5753 ( .D(g2142), .ISO(n3425), .Q(n3424) );
  ISOLANDX1 U5754 ( .D(g2151), .ISO(n3684), .Q(n3683) );
  ISOLANDX1 U5755 ( .D(g2160), .ISO(n3888), .Q(n3887) );
  ISOLANDX1 U5756 ( .D(g1448), .ISO(n3428), .Q(n3427) );
  ISOLANDX1 U5757 ( .D(g1457), .ISO(n3687), .Q(n3686) );
  ISOLANDX1 U5758 ( .D(g1466), .ISO(n3891), .Q(n3890) );
  ISOLANDX1 U5759 ( .D(g762), .ISO(n3431), .Q(n3430) );
  ISOLANDX1 U5760 ( .D(g771), .ISO(n3690), .Q(n3689) );
  ISOLANDX1 U5761 ( .D(g780), .ISO(n3894), .Q(n3893) );
  ISOLANDX1 U5762 ( .D(g74), .ISO(n3434), .Q(n3433) );
  ISOLANDX1 U5763 ( .D(g83), .ISO(n3693), .Q(n3692) );
  ISOLANDX1 U5764 ( .D(g92), .ISO(n3897), .Q(n3896) );
  NOR2X0 U5765 ( .IN1(n3739), .IN2(n3740), .QN(g26786) );
  XOR2X1 U5766 ( .IN1(n3741), .IN2(g3024), .Q(n3739) );
  NOR2X0 U5767 ( .IN1(n3861), .IN2(n3740), .QN(g26031) );
  XOR2X1 U5768 ( .IN1(n3742), .IN2(test_so98), .Q(n3861) );
  NOR2X0 U5769 ( .IN1(n4103), .IN2(n3740), .QN(g24445) );
  XOR2X1 U5770 ( .IN1(n4066), .IN2(g3002), .Q(n4103) );
  NAND4X0 U5771 ( .IN1(n4305), .IN2(n4355), .IN3(n4291), .IN4(n4223), .QN(
        n2505) );
  NAND2X0 U5772 ( .IN1(n3858), .IN2(n3994), .QN(g25265) );
  NAND3X0 U5773 ( .IN1(n3995), .IN2(n3859), .IN3(n1581), .QN(n3994) );
  OR2X1 U5774 ( .IN1(g2993), .IN2(n4597), .Q(n3995) );
  OA22X1_S38584 U5775 ( .IN1(n2487), .IN2(n2488), .IN3(n2489), .IN4(n2490), .Q(n4275)
         );
  NAND4X0 U5776 ( .IN1(n2504), .IN2(n4651), .IN3(n2506), .IN4(n2507), .QN(
        n2487) );
  NAND4X0 U5777 ( .IN1(n2491), .IN2(n2492), .IN3(n2493), .IN4(n2494), .QN(
        n2488) );
  XOR2X1 U5778 ( .IN1(g2147), .IN2(n2078), .Q(n2506) );
  OA22X1_S38584 U5779 ( .IN1(n2514), .IN2(n2515), .IN3(n2516), .IN4(n2517), .Q(n4276)
         );
  NAND4X0 U5780 ( .IN1(n2531), .IN2(n4651), .IN3(n2532), .IN4(n2533), .QN(
        n2514) );
  NAND4X0 U5781 ( .IN1(n2518), .IN2(n2519), .IN3(n2520), .IN4(n2521), .QN(
        n2515) );
  XOR2X1 U5782 ( .IN1(g1453), .IN2(n1976), .Q(n2532) );
  OA22X1_S38584 U5783 ( .IN1(n2540), .IN2(n2541), .IN3(n2542), .IN4(n2543), .Q(n4277)
         );
  NAND4X0 U5784 ( .IN1(n2557), .IN2(n4651), .IN3(n2558), .IN4(n2559), .QN(
        n2540) );
  NAND4X0 U5785 ( .IN1(n2544), .IN2(n2545), .IN3(n2546), .IN4(n2547), .QN(
        n2541) );
  XOR2X1 U5786 ( .IN1(g767), .IN2(n1875), .Q(n2558) );
  OA22X1_S38584 U5787 ( .IN1(n2566), .IN2(n2567), .IN3(n2568), .IN4(n2569), .Q(n4278)
         );
  NAND4X0 U5788 ( .IN1(n2583), .IN2(n4651), .IN3(n2584), .IN4(n2585), .QN(
        n2566) );
  NAND4X0 U5789 ( .IN1(n2570), .IN2(n2571), .IN3(n2572), .IN4(n2573), .QN(
        n2567) );
  XOR2X1 U5790 ( .IN1(test_so15), .IN2(n1770), .Q(n2584) );
  OA22X1_S38584 U5791 ( .IN1(g2652), .IN2(n2122), .IN3(n3511), .IN4(n3503), .Q(g27343) );
  OA22X1_S38584 U5792 ( .IN1(g2654), .IN2(n2123), .IN3(n3511), .IN4(n3504), .Q(g27337) );
  OA22X1_S38584 U5793 ( .IN1(g2653), .IN2(n2121), .IN3(n3511), .IN4(n3508), .Q(g27326) );
  OA22X1_S38584 U5794 ( .IN1(g1958), .IN2(n2020), .IN3(n3528), .IN4(n3507), .Q(g27331) );
  OA22X1_S38584 U5795 ( .IN1(g1960), .IN2(n2021), .IN3(n3528), .IN4(n3514), .Q(g27320) );
  OA22X1_S38584 U5796 ( .IN1(g1959), .IN2(n2019), .IN3(n3528), .IN4(n3525), .Q(g27306) );
  OA22X1_S38584 U5797 ( .IN1(g1264), .IN2(n1918), .IN3(n3554), .IN4(n3517), .Q(g27314) );
  OA22X1_S38584 U5798 ( .IN1(g1266), .IN2(n1919), .IN3(n3554), .IN4(n3531), .Q(g27300) );
  OA22X1_S38584 U5799 ( .IN1(g1265), .IN2(n1917), .IN3(n3554), .IN4(n3551), .Q(g27286) );
  OA22X1_S38584 U5800 ( .IN1(g578), .IN2(n1814), .IN3(n3589), .IN4(n3534), .Q(g27294)
         );
  OA22X1_S38584 U5801 ( .IN1(test_so25), .IN2(n1815), .IN3(n3589), .IN4(n3557), .Q(
        g27280) );
  OA22X1_S38584 U5802 ( .IN1(g579), .IN2(n1813), .IN3(n3589), .IN4(n3586), .Q(g27269)
         );
  OA22X1_S38584 U5803 ( .IN1(g2658), .IN2(n2122), .IN3(n3502), .IN4(n3503), .Q(g27354) );
  OA22X1_S38584 U5804 ( .IN1(g2660), .IN2(n2123), .IN3(n3502), .IN4(n3504), .Q(g27348) );
  OA22X1_S38584 U5805 ( .IN1(g2659), .IN2(n2121), .IN3(n3502), .IN4(n3508), .Q(g27345) );
  OA22X1_S38584 U5806 ( .IN1(g1964), .IN2(n2020), .IN3(n3506), .IN4(n3507), .Q(g27346) );
  OA22X1_S38584 U5807 ( .IN1(g1966), .IN2(n2021), .IN3(n3506), .IN4(n3514), .Q(g27341) );
  OA22X1_S38584 U5808 ( .IN1(test_so67), .IN2(n2019), .IN3(n3506), .IN4(n3525), .Q(
        g27333) );
  OA22X1_S38584 U5809 ( .IN1(g1270), .IN2(n1918), .IN3(n3516), .IN4(n3517), .Q(g27339) );
  OA22X1_S38584 U5810 ( .IN1(g1272), .IN2(n1919), .IN3(n3516), .IN4(n3531), .Q(g27329) );
  OA22X1_S38584 U5811 ( .IN1(g1271), .IN2(n1917), .IN3(n3516), .IN4(n3551), .Q(g27316) );
  OA22X1_S38584 U5812 ( .IN1(g584), .IN2(n1814), .IN3(n3533), .IN4(n3534), .Q(g27327)
         );
  OA22X1_S38584 U5813 ( .IN1(g586), .IN2(n1815), .IN3(n3533), .IN4(n3557), .Q(g27312)
         );
  OA22X1_S38584 U5814 ( .IN1(g585), .IN2(n1813), .IN3(n3533), .IN4(n3586), .Q(g27296)
         );
  OA22X1_S38584 U5815 ( .IN1(g2655), .IN2(n2122), .IN3(n3505), .IN4(n3503), .Q(g27347) );
  OA22X1_S38584 U5816 ( .IN1(test_so89), .IN2(n2123), .IN3(n3505), .IN4(n3504), .Q(
        g27344) );
  OA22X1_S38584 U5817 ( .IN1(g2656), .IN2(n2121), .IN3(n3505), .IN4(n3508), .Q(g27338) );
  OA22X1_S38584 U5818 ( .IN1(g2649), .IN2(n2122), .IN3(n3522), .IN4(n3503), .Q(g27336) );
  OA22X1_S38584 U5819 ( .IN1(g2651), .IN2(n2123), .IN3(n3522), .IN4(n3504), .Q(g27325) );
  OA22X1_S38584 U5820 ( .IN1(g2650), .IN2(n2121), .IN3(n3522), .IN4(n3508), .Q(g27310) );
  OA22X1_S38584 U5821 ( .IN1(g1961), .IN2(n2020), .IN3(n3515), .IN4(n3507), .Q(g27340) );
  OA22X1_S38584 U5822 ( .IN1(g1963), .IN2(n2021), .IN3(n3515), .IN4(n3514), .Q(g27332) );
  OA22X1_S38584 U5823 ( .IN1(g1962), .IN2(n2019), .IN3(n3515), .IN4(n3525), .Q(g27321) );
  OA22X1_S38584 U5824 ( .IN1(g1955), .IN2(n2020), .IN3(n3548), .IN4(n3507), .Q(g27319) );
  OA22X1_S38584 U5825 ( .IN1(g1957), .IN2(n2021), .IN3(n3548), .IN4(n3514), .Q(g27305) );
  OA22X1_S38584 U5826 ( .IN1(g1956), .IN2(n2019), .IN3(n3548), .IN4(n3525), .Q(g27290) );
  OA22X1_S38584 U5827 ( .IN1(test_so46), .IN2(n1918), .IN3(n3532), .IN4(n3517), .Q(
        g27328) );
  OA22X1_S38584 U5828 ( .IN1(g1269), .IN2(n1919), .IN3(n3532), .IN4(n3531), .Q(g27315) );
  OA22X1_S38584 U5829 ( .IN1(g1268), .IN2(n1917), .IN3(n3532), .IN4(n3551), .Q(g27301) );
  OA22X1_S38584 U5830 ( .IN1(g1261), .IN2(n1918), .IN3(n3583), .IN4(n3517), .Q(g27299) );
  OA22X1_S38584 U5831 ( .IN1(g1263), .IN2(n1919), .IN3(n3583), .IN4(n3531), .Q(g27285) );
  OA22X1_S38584 U5832 ( .IN1(g1262), .IN2(n1917), .IN3(n3583), .IN4(n3551), .Q(g27273) );
  OA22X1_S38584 U5833 ( .IN1(g581), .IN2(n1814), .IN3(n3558), .IN4(n3534), .Q(g27311)
         );
  OA22X1_S38584 U5834 ( .IN1(g583), .IN2(n1815), .IN3(n3558), .IN4(n3557), .Q(g27295)
         );
  OA22X1_S38584 U5835 ( .IN1(g582), .IN2(n1813), .IN3(n3558), .IN4(n3586), .Q(g27281)
         );
  OA22X1_S38584 U5836 ( .IN1(g575), .IN2(n1814), .IN3(n3619), .IN4(n3534), .Q(g27279)
         );
  OA22X1_S38584 U5837 ( .IN1(g577), .IN2(n1815), .IN3(n3619), .IN4(n3557), .Q(g27268)
         );
  OA22X1_S38584 U5838 ( .IN1(g576), .IN2(n1813), .IN3(n3619), .IN4(n3586), .Q(g27261)
         );
  OA21X1 U5839 ( .IN1(n4306), .IN2(g2809), .IN3(n2388), .Q(n2387) );
  OA21X1 U5840 ( .IN1(n4307), .IN2(g2115), .IN3(n2316), .Q(n2315) );
  OA21X1 U5841 ( .IN1(n4308), .IN2(g1421), .IN3(n2244), .Q(n2243) );
  OA21X1 U5842 ( .IN1(n4309), .IN2(g735), .IN3(n2451), .Q(n2450) );
  OAI222X1 U5843 ( .IN1(n4359), .IN2(g739), .IN3(n4309), .IN4(g738), .IN5(
        n4295), .IN6(g737), .QN(n2477) );
  OAI222X1 U5844 ( .IN1(n4356), .IN2(g2813), .IN3(n4306), .IN4(g2812), .IN5(
        n4292), .IN6(test_so95), .QN(n2399) );
  OAI222X1 U5845 ( .IN1(n4357), .IN2(g2119), .IN3(n4307), .IN4(g2118), .IN5(
        n4293), .IN6(g2117), .QN(n2327) );
  OAI222X1 U5846 ( .IN1(n4358), .IN2(g1425), .IN3(n4308), .IN4(g1424), .IN5(
        n4294), .IN6(g1423), .QN(n2255) );
  NOR3X0 U5847 ( .IN1(n2548), .IN2(n2549), .IN3(n2550), .QN(n2547) );
  XNOR2X1 U5848 ( .IN1(n2552), .IN2(g740), .Q(n2549) );
  XOR2X1 U5849 ( .IN1(n2551), .IN2(g771), .Q(n2550) );
  XNOR2X1 U5850 ( .IN1(n2553), .IN2(g744), .Q(n2548) );
  NBUFFX2 U5851 ( .IN(g2480), .Q(g7264) );
  NBUFFX2 U5852 ( .IN(g1786), .Q(g7014) );
  NBUFFX2 U5853 ( .IN(g2351), .Q(g5555) );
  NBUFFX2 U5854 ( .IN(g1657), .Q(g5511) );
  NBUFFX2 U5855 ( .IN(g276), .Q(g5437) );
  NBUFFX2 U5856 ( .IN(g1925), .Q(n4616) );
  NBUFFX2 U5857 ( .IN(g1231), .Q(n4628) );
  AO222X1 U5858 ( .IN1(g2584), .IN2(n2329), .IN3(n2330), .IN4(n1570), .IN5(
        g2631), .IN6(n2331), .Q(n4250) );
  NOR2X0 U5859 ( .IN1(n2137), .IN2(n2334), .QN(n2330) );
  XOR2X1 U5860 ( .IN1(n2332), .IN2(n2333), .Q(n2331) );
  XOR2X1 U5861 ( .IN1(n2335), .IN2(n2336), .Q(n2329) );
  AO222X1 U5862 ( .IN1(g1890), .IN2(n2257), .IN3(n2258), .IN4(n1568), .IN5(
        g1937), .IN6(n2259), .Q(n4241) );
  NOR2X0 U5863 ( .IN1(n2035), .IN2(n2262), .QN(n2258) );
  XOR2X1 U5864 ( .IN1(n2260), .IN2(n2261), .Q(n2259) );
  XOR2X1 U5865 ( .IN1(n2263), .IN2(n2264), .Q(n2257) );
  NOR3X0 U5866 ( .IN1(n2495), .IN2(n2496), .IN3(n2497), .QN(n2494) );
  XNOR2X1 U5867 ( .IN1(n2499), .IN2(g2120), .Q(n2496) );
  XOR2X1 U5868 ( .IN1(n2498), .IN2(g2151), .Q(n2497) );
  XOR2X1 U5869 ( .IN1(n2500), .IN2(g2124), .Q(n2495) );
  NOR3X0 U5870 ( .IN1(n2522), .IN2(n2523), .IN3(n2524), .QN(n2521) );
  XNOR2X1 U5871 ( .IN1(n2526), .IN2(g1426), .Q(n2523) );
  XOR2X1 U5872 ( .IN1(n2525), .IN2(g1457), .Q(n2524) );
  XOR2X1 U5873 ( .IN1(n2527), .IN2(g1430), .Q(n2522) );
  NOR3X0 U5874 ( .IN1(n2574), .IN2(n2575), .IN3(n2576), .QN(n2573) );
  XNOR2X1 U5875 ( .IN1(n2578), .IN2(g52), .Q(n2575) );
  XOR2X1 U5876 ( .IN1(n2577), .IN2(g83), .Q(n2576) );
  XOR2X1 U5877 ( .IN1(n2579), .IN2(g56), .Q(n2574) );
  NBUFFX2 U5878 ( .IN(g2476), .Q(n4605) );
  NBUFFX2 U5879 ( .IN(g1782), .Q(n4617) );
  NBUFFX2 U5880 ( .IN(g401), .Q(n4639) );
  NOR3X0 U5881 ( .IN1(n4056), .IN2(n1580), .IN3(n4101), .QN(g24446) );
  ISOLANDX1 U5882 ( .D(n4102), .ISO(g3036), .Q(n4101) );
  NOR2X0 U5883 ( .IN1(n1580), .IN2(n4055), .QN(g25202) );
  XNOR2X1 U5884 ( .IN1(g3032), .IN2(n4056), .Q(n4055) );
  NOR2X0 U5885 ( .IN1(n1606), .IN2(n2980), .QN(g29582) );
  XOR2X1 U5886 ( .IN1(n2981), .IN2(g2120), .Q(n2980) );
  NOR2X0 U5887 ( .IN1(n1605), .IN2(n2983), .QN(g29581) );
  XOR2X1 U5888 ( .IN1(n2984), .IN2(g1426), .Q(n2983) );
  NOR2X0 U5889 ( .IN1(n1604), .IN2(n2986), .QN(g29580) );
  XOR2X1 U5890 ( .IN1(n2987), .IN2(g740), .Q(n2986) );
  NOR2X0 U5891 ( .IN1(n1603), .IN2(n2989), .QN(g29579) );
  XOR2X1 U5892 ( .IN1(n2990), .IN2(g52), .Q(n2989) );
  OA222X1 U5893 ( .IN1(n4370), .IN2(test_so89), .IN3(n4299), .IN4(g2655), 
        .IN5(n4314), .IN6(g2656), .Q(n3279) );
  OA222X1 U5894 ( .IN1(n4315), .IN2(g1963), .IN3(n4366), .IN4(g1961), .IN5(
        n4296), .IN6(g1962), .Q(n3320) );
  OA222X1 U5895 ( .IN1(n4316), .IN2(g1269), .IN3(n4300), .IN4(test_so46), 
        .IN5(n4371), .IN6(g1268), .Q(n3360) );
  OA222X1 U5896 ( .IN1(n4372), .IN2(g583), .IN3(n4313), .IN4(g581), .IN5(n4298), .IN6(g582), .Q(n3399) );
  AO222X1 U5897 ( .IN1(g2441), .IN2(g5796), .IN3(g2443), .IN4(g2412), .IN5(
        g2439), .IN6(g5747), .Q(n3277) );
  AO222X1 U5898 ( .IN1(g1747), .IN2(g5738), .IN3(g1749), .IN4(g1718), .IN5(
        g1745), .IN6(g5695), .Q(n3318) );
  AO222X1 U5899 ( .IN1(g1053), .IN2(g5686), .IN3(g1055), .IN4(g1024), .IN5(
        g1051), .IN6(g5657), .Q(n3358) );
  AO222X1 U5900 ( .IN1(g366), .IN2(g5648), .IN3(g368), .IN4(g337), .IN5(g364), 
        .IN6(g5629), .Q(n3397) );
  OA222X1 U5901 ( .IN1(n4673), .IN2(g1002), .IN3(n4669), .IN4(g1004), .IN5(
        n4671), .IN6(g1003), .Q(n2618) );
  OA222X1 U5902 ( .IN1(n4673), .IN2(g1005), .IN3(n4669), .IN4(test_so39), 
        .IN5(n4671), .IN6(g1006), .Q(n2627) );
  OA222X1 U5903 ( .IN1(n4682), .IN2(g2252), .IN3(n4680), .IN4(g2250), .IN5(
        n4683), .IN6(g2251), .Q(n3062) );
  OA222X1 U5904 ( .IN1(n4686), .IN2(g1558), .IN3(n4685), .IN4(g1556), .IN5(
        n4317), .IN6(g1557), .Q(n3094) );
  OA222X1 U5905 ( .IN1(n4696), .IN2(g176), .IN3(n4695), .IN4(g174), .IN5(n4318), .IN6(g175), .Q(n3154) );
  OA222X1 U5906 ( .IN1(n4312), .IN2(g864), .IN3(n4362), .IN4(g862), .IN5(n4693), .IN6(g863), .Q(n3227) );
  OA222X1 U5907 ( .IN1(n4673), .IN2(g999), .IN3(n4669), .IN4(g1001), .IN5(
        n4671), .IN6(g1000), .Q(n4118) );
  AO222X1 U5908 ( .IN1(g921), .IN2(n4591), .IN3(test_so34), .IN4(test_so31), 
        .IN5(g918), .IN6(n4592), .Q(n2564) );
  AO222X1 U5909 ( .IN1(g930), .IN2(n4591), .IN3(g933), .IN4(test_so31), .IN5(
        g927), .IN6(n4592), .Q(n2743) );
  AO222X1 U5910 ( .IN1(g2471), .IN2(g5796), .IN3(test_so85), .IN4(g2412), 
        .IN5(g2469), .IN6(g5747), .Q(n3270) );
  OA222X1 U5911 ( .IN1(n4664), .IN2(g2398), .IN3(n4663), .IN4(g2396), .IN5(
        n4665), .IN6(g2397), .Q(n2898) );
  OA222X1 U5912 ( .IN1(n4667), .IN2(g1704), .IN3(n4666), .IN4(g1702), .IN5(
        n4668), .IN6(g1703), .Q(n2916) );
  OA222X1 U5913 ( .IN1(n4674), .IN2(g1009), .IN3(n4670), .IN4(g1008), .IN5(
        n4672), .IN6(g1010), .Q(n2934) );
  OA222X1 U5914 ( .IN1(n4677), .IN2(g323), .IN3(n4675), .IN4(g321), .IN5(n4678), .IN6(g322), .Q(n2951) );
  AO222X1 U5915 ( .IN1(g885), .IN2(g6518), .IN3(g888), .IN4(test_so31), .IN5(
        g882), .IN6(g6368), .Q(n2551) );
  AO222X1 U5916 ( .IN1(g876), .IN2(n4591), .IN3(g879), .IN4(n4689), .IN5(g873), 
        .IN6(n4592), .Q(n2565) );
  OA222X1 U5917 ( .IN1(n4682), .IN2(g2249), .IN3(n4680), .IN4(g2247), .IN5(
        n4683), .IN6(g2248), .Q(n2666) );
  OA222X1 U5918 ( .IN1(n4686), .IN2(g1555), .IN3(n4685), .IN4(test_so54), 
        .IN5(n4317), .IN6(g1554), .Q(n2681) );
  OA222X1 U5919 ( .IN1(n4312), .IN2(g861), .IN3(n4362), .IN4(g859), .IN5(n4693), .IN6(g860), .Q(n2696) );
  OA222X1 U5920 ( .IN1(n4696), .IN2(g173), .IN3(n4695), .IN4(g171), .IN5(n4318), .IN6(g172), .Q(n2714) );
  XOR2X1 U5921 ( .IN1(n2511), .IN2(g2185), .Q(n3043) );
  XOR2X1 U5922 ( .IN1(n2537), .IN2(g1491), .Q(n3075) );
  XOR2X1 U5923 ( .IN1(n2563), .IN2(g801), .Q(n3107) );
  XOR2X1 U5924 ( .IN1(n2589), .IN2(g113), .Q(n3135) );
  AO222X1 U5925 ( .IN1(g903), .IN2(n4591), .IN3(g906), .IN4(n4689), .IN5(g900), 
        .IN6(n4592), .Q(n2554) );
  AO222X1 U5926 ( .IN1(g948), .IN2(n4591), .IN3(g951), .IN4(n4689), .IN5(
        test_so35), .IN6(n4592), .Q(n2555) );
  AO222X1 U5927 ( .IN1(g939), .IN2(g6518), .IN3(g942), .IN4(test_so31), .IN5(
        g936), .IN6(g6368), .Q(n2556) );
  XOR2X1 U5928 ( .IN1(n2503), .IN2(g2190), .Q(n3060) );
  XOR2X1 U5929 ( .IN1(n2530), .IN2(g1496), .Q(n3092) );
  XOR2X1 U5930 ( .IN1(n2556), .IN2(g805), .Q(n3124) );
  XOR2X1 U5931 ( .IN1(n2582), .IN2(g117), .Q(n3152) );
  INVX0 U5932 ( .IN(test_so31), .QN(n4691) );
  OA222X1 U5933 ( .IN1(n4681), .IN2(g2246), .IN3(n4680), .IN4(g2244), .IN5(
        n4683), .IN6(g2245), .Q(n3199) );
  OA222X1 U5934 ( .IN1(n4686), .IN2(g1552), .IN3(n4685), .IN4(g1550), .IN5(
        n4317), .IN6(g1551), .Q(n3215) );
  OA222X1 U5935 ( .IN1(n4312), .IN2(test_so33), .IN3(n4362), .IN4(g856), .IN5(
        n4693), .IN6(g857), .Q(n3229) );
  OA222X1 U5936 ( .IN1(n4696), .IN2(g170), .IN3(n4695), .IN4(g168), .IN5(n4318), .IN6(g169), .Q(n3240) );
  AOI222X1 U5937 ( .IN1(g912), .IN2(g6518), .IN3(g915), .IN4(n4689), .IN5(g909), .IN6(g6368), .QN(n2553) );
  AOI222X1 U5938 ( .IN1(g894), .IN2(g6518), .IN3(g897), .IN4(n4689), .IN5(g891), .IN6(g6368), .QN(n2563) );
  ISOLANDX1 U5939 ( .D(g2257), .ISO(n3199), .Q(n3038) );
  ISOLANDX1 U5940 ( .D(g1563), .ISO(n3215), .Q(n3070) );
  ISOLANDX1 U5941 ( .D(g869), .ISO(n3229), .Q(n3102) );
  ISOLANDX1 U5942 ( .D(g181), .ISO(n3240), .Q(n3130) );
  AO221X1 U5943 ( .IN1(n2659), .IN2(g2175), .IN3(n2660), .IN4(n2661), .IN5(
        n2662), .Q(n2656) );
  XOR2X1 U5944 ( .IN1(n2663), .IN2(n2498), .Q(n2660) );
  AO221X1 U5945 ( .IN1(n2673), .IN2(g1481), .IN3(n2674), .IN4(n2675), .IN5(
        n2676), .Q(n2658) );
  XOR2X1 U5946 ( .IN1(n2677), .IN2(n2525), .Q(n2674) );
  AO221X1 U5947 ( .IN1(n2688), .IN2(g793), .IN3(n2689), .IN4(n2690), .IN5(
        n2691), .Q(n2665) );
  XOR2X1 U5948 ( .IN1(n2692), .IN2(n2551), .Q(n2689) );
  AO221X1 U5949 ( .IN1(n2702), .IN2(g105), .IN3(n2703), .IN4(n2704), .IN5(
        n2705), .Q(n2679) );
  XOR2X1 U5950 ( .IN1(n2706), .IN2(n2577), .Q(n2703) );
  OA222X1 U5951 ( .IN1(g2235), .IN2(n4680), .IN3(g2237), .IN4(n4681), .IN5(
        g2236), .IN6(n4683), .Q(n3885) );
  OA222X1 U5952 ( .IN1(g1541), .IN2(n4685), .IN3(g1543), .IN4(n4686), .IN5(
        g1542), .IN6(n4317), .Q(n3782) );
  OA222X1 U5953 ( .IN1(g847), .IN2(n4362), .IN3(g849), .IN4(n4692), .IN5(g848), 
        .IN6(n4693), .Q(n3812) );
  OA222X1 U5954 ( .IN1(g159), .IN2(n4695), .IN3(g161), .IN4(n4696), .IN5(g160), 
        .IN6(n4318), .Q(n3840) );
  OA222X1 U5955 ( .IN1(g2238), .IN2(n4680), .IN3(test_so75), .IN4(n4681), 
        .IN5(g2239), .IN6(n4324), .Q(n3884) );
  OA222X1 U5956 ( .IN1(g1544), .IN2(n4685), .IN3(g1546), .IN4(n4686), .IN5(
        g1545), .IN6(n4688), .Q(n3781) );
  OA222X1 U5957 ( .IN1(g850), .IN2(n4362), .IN3(g852), .IN4(n4312), .IN5(g851), 
        .IN6(n4323), .Q(n3811) );
  OA222X1 U5958 ( .IN1(g162), .IN2(n4695), .IN3(g164), .IN4(n4696), .IN5(
        test_so12), .IN6(n4698), .Q(n3839) );
  AO22X1 U5959 ( .IN1(n2890), .IN2(n2661), .IN3(n2659), .IN4(g2195), .Q(n2880)
         );
  XOR2X1 U5960 ( .IN1(n2736), .IN2(n2501), .Q(n2890) );
  AO22X1 U5961 ( .IN1(n2842), .IN2(n2661), .IN3(n2659), .IN4(g2185), .Q(n2840)
         );
  XNOR2X1 U5962 ( .IN1(n2511), .IN2(n2843), .Q(n2842) );
  AO22X1 U5963 ( .IN1(n2908), .IN2(n2675), .IN3(n2673), .IN4(g1501), .Q(n2886)
         );
  XOR2X1 U5964 ( .IN1(n2751), .IN2(n2528), .Q(n2908) );
  AO22X1 U5965 ( .IN1(n2847), .IN2(n2675), .IN3(n2673), .IN4(g1491), .Q(n2841)
         );
  XNOR2X1 U5966 ( .IN1(n2537), .IN2(n2848), .Q(n2847) );
  AO22X1 U5967 ( .IN1(n2926), .IN2(n2690), .IN3(n2688), .IN4(g809), .Q(n2907)
         );
  XOR2X1 U5968 ( .IN1(n2766), .IN2(n2554), .Q(n2926) );
  AO22X1 U5969 ( .IN1(n2854), .IN2(n2690), .IN3(n2688), .IN4(g801), .Q(n2845)
         );
  XNOR2X1 U5970 ( .IN1(n2563), .IN2(n2855), .Q(n2854) );
  AO22X1 U5971 ( .IN1(n2943), .IN2(n2704), .IN3(n2702), .IN4(g121), .Q(n2925)
         );
  XOR2X1 U5972 ( .IN1(n2775), .IN2(n2580), .Q(n2943) );
  AO22X1 U5973 ( .IN1(n2862), .IN2(n2704), .IN3(n2702), .IN4(g113), .Q(n2850)
         );
  XNOR2X1 U5974 ( .IN1(n2589), .IN2(n2863), .Q(n2862) );
  AO22X1 U5975 ( .IN1(n2661), .IN2(n2852), .IN3(n2659), .IN4(g2165), .Q(n2844)
         );
  XOR2X1 U5976 ( .IN1(n2513), .IN2(n2725), .Q(n2852) );
  AO22X1 U5977 ( .IN1(n2675), .IN2(n2860), .IN3(n2673), .IN4(g1471), .Q(n2849)
         );
  XOR2X1 U5978 ( .IN1(n2539), .IN2(n2741), .Q(n2860) );
  AO22X1 U5979 ( .IN1(n2690), .IN2(n2871), .IN3(n2688), .IN4(g785), .Q(n2856)
         );
  XOR2X1 U5980 ( .IN1(n2565), .IN2(n2757), .Q(n2871) );
  AO22X1 U5981 ( .IN1(n2704), .IN2(n2879), .IN3(n2702), .IN4(g97), .Q(n2864)
         );
  XOR2X1 U5982 ( .IN1(n2591), .IN2(n2771), .Q(n2879) );
  AOI222X1 U5983 ( .IN1(g1651), .IN2(n4589), .IN3(g1654), .IN4(n4684), .IN5(
        g1648), .IN6(g6573), .QN(n2526) );
  AOI222X1 U5984 ( .IN1(g957), .IN2(n4591), .IN3(g960), .IN4(n4689), .IN5(g954), .IN6(n4592), .QN(n2552) );
  AOI222X1 U5985 ( .IN1(g270), .IN2(n4593), .IN3(g273), .IN4(n4694), .IN5(g267), .IN6(g6231), .QN(n2578) );
  XOR2X1 U5986 ( .IN1(n2076), .IN2(g2170), .Q(n3057) );
  XOR2X1 U5987 ( .IN1(n1974), .IN2(g1476), .Q(n3089) );
  XOR2X1 U5988 ( .IN1(n1873), .IN2(g789), .Q(n3121) );
  XOR2X1 U5989 ( .IN1(n1768), .IN2(g101), .Q(n3149) );
  XOR2X1 U5990 ( .IN1(n2078), .IN2(g2180), .Q(n3054) );
  XOR2X1 U5991 ( .IN1(n1976), .IN2(g1486), .Q(n3086) );
  XOR2X1 U5992 ( .IN1(n2079), .IN2(g2175), .Q(n3044) );
  XOR2X1 U5993 ( .IN1(n1977), .IN2(g1481), .Q(n3076) );
  XOR2X1 U5994 ( .IN1(n1875), .IN2(g797), .Q(n3118) );
  XOR2X1 U5995 ( .IN1(n1770), .IN2(g109), .Q(n3146) );
  XOR2X1 U5996 ( .IN1(n1876), .IN2(g793), .Q(n3108) );
  XOR2X1 U5997 ( .IN1(n1771), .IN2(g105), .Q(n3136) );
  XOR2X1 U5998 ( .IN1(n2077), .IN2(g2165), .Q(n3047) );
  XOR2X1 U5999 ( .IN1(n1975), .IN2(g1471), .Q(n3079) );
  XOR2X1 U6000 ( .IN1(n1874), .IN2(g785), .Q(n3111) );
  XOR2X1 U6001 ( .IN1(n4513), .IN2(g97), .Q(n3139) );
  AO22X1 U6002 ( .IN1(g2330), .IN2(n4367), .IN3(n2851), .IN4(g2241), .Q(g30290) );
  AO22X1 U6003 ( .IN1(g2321), .IN2(n4680), .IN3(n2680), .IN4(g2241), .Q(g30679) );
  AO22X1 U6004 ( .IN1(g2312), .IN2(n4680), .IN3(n2694), .IN4(g2241), .Q(g30672) );
  AO22X1 U6005 ( .IN1(g1636), .IN2(n4368), .IN3(n2859), .IN4(g1547), .Q(g30280) );
  AO22X1 U6006 ( .IN1(g1627), .IN2(n4685), .IN3(n2695), .IN4(g1547), .Q(g30671) );
  AO22X1 U6007 ( .IN1(g1618), .IN2(n4685), .IN3(n2712), .IN4(g1547), .Q(g30663) );
  AO22X1 U6008 ( .IN1(g960), .IN2(n4362), .IN3(n2678), .IN4(n4690), .Q(g30682)
         );
  AO22X1 U6009 ( .IN1(g951), .IN2(n4691), .IN3(n2861), .IN4(n4690), .Q(g30278)
         );
  AO22X1 U6010 ( .IN1(g942), .IN2(n4691), .IN3(n2870), .IN4(n4690), .Q(g30270)
         );
  AO22X1 U6011 ( .IN1(g933), .IN2(n4362), .IN3(n2713), .IN4(n4690), .Q(g30662)
         );
  AO22X1 U6012 ( .IN1(test_so34), .IN2(n4362), .IN3(n2731), .IN4(n4690), .Q(
        g30654) );
  AO22X1 U6013 ( .IN1(test_so14), .IN2(n4369), .IN3(n2878), .IN4(g165), .Q(
        g30262) );
  AO22X1 U6014 ( .IN1(g246), .IN2(n4695), .IN3(n2732), .IN4(g165), .Q(g30653)
         );
  AO22X1 U6015 ( .IN1(g237), .IN2(n4695), .IN3(n2747), .IN4(g165), .Q(g30645)
         );
  AO22X1 U6016 ( .IN1(g2336), .IN2(n4681), .IN3(n2846), .IN4(n4587), .Q(g30291) );
  AO22X1 U6017 ( .IN1(g2333), .IN2(n4324), .IN3(n2846), .IN4(g6837), .Q(g30283) );
  AO22X1 U6018 ( .IN1(g2291), .IN2(n4681), .IN3(g7084), .IN4(n2880), .Q(g30256) );
  AO22X1 U6019 ( .IN1(g2288), .IN2(n4324), .IN3(g2214), .IN4(n2880), .Q(g30253) );
  AO22X1 U6020 ( .IN1(test_so77), .IN2(n4681), .IN3(n2851), .IN4(g7084), .Q(
        g30282) );
  AO22X1 U6021 ( .IN1(g2324), .IN2(n4324), .IN3(n2851), .IN4(g2214), .Q(g30274) );
  AO22X1 U6022 ( .IN1(g2282), .IN2(n4681), .IN3(n4587), .IN4(n2840), .Q(g30303) );
  AO22X1 U6023 ( .IN1(g2279), .IN2(n4683), .IN3(g6837), .IN4(n2840), .Q(g30301) );
  AO22X1 U6024 ( .IN1(g2315), .IN2(n4683), .IN3(n2680), .IN4(g6837), .Q(g30667) );
  AO22X1 U6025 ( .IN1(g2273), .IN2(n4681), .IN3(g7084), .IN4(n2656), .Q(g30693) );
  AO22X1 U6026 ( .IN1(g2270), .IN2(n4324), .IN3(g2214), .IN4(n2656), .Q(g30690) );
  AO22X1 U6027 ( .IN1(g2306), .IN2(n4683), .IN3(n2694), .IN4(g6837), .Q(g30660) );
  AO22X1 U6028 ( .IN1(test_so76), .IN2(n4681), .IN3(n4587), .IN4(n2844), .Q(
        g30296) );
  AO22X1 U6029 ( .IN1(g2261), .IN2(n4683), .IN3(g2214), .IN4(n2844), .Q(g30289) );
  AO22X1 U6030 ( .IN1(g1642), .IN2(n4687), .IN3(n2853), .IN4(n4589), .Q(g30281) );
  AO22X1 U6031 ( .IN1(g1639), .IN2(n4688), .IN3(n2853), .IN4(g6573), .Q(g30273) );
  AO22X1 U6032 ( .IN1(g1597), .IN2(n4687), .IN3(g6782), .IN4(n2886), .Q(g30252) );
  AO22X1 U6033 ( .IN1(g1594), .IN2(n4688), .IN3(g1520), .IN4(n2886), .Q(g30250) );
  AO22X1 U6034 ( .IN1(g1633), .IN2(n4687), .IN3(n2859), .IN4(g6782), .Q(g30272) );
  AO22X1 U6035 ( .IN1(g1630), .IN2(n4688), .IN3(n2859), .IN4(g1520), .Q(g30266) );
  AO22X1 U6036 ( .IN1(g1588), .IN2(n4687), .IN3(n4589), .IN4(n2841), .Q(g30299) );
  AO22X1 U6037 ( .IN1(g1585), .IN2(n4317), .IN3(g6573), .IN4(n2841), .Q(g30295) );
  AO22X1 U6038 ( .IN1(test_so55), .IN2(n4317), .IN3(n2695), .IN4(g6573), .Q(
        g30658) );
  AO22X1 U6039 ( .IN1(g1579), .IN2(n4687), .IN3(n4589), .IN4(n2658), .Q(g30688) );
  AO22X1 U6040 ( .IN1(g1576), .IN2(n4688), .IN3(g1520), .IN4(n2658), .Q(g30683) );
  AO22X1 U6041 ( .IN1(g1612), .IN2(n4317), .IN3(n2712), .IN4(g6573), .Q(g30651) );
  AO22X1 U6042 ( .IN1(g1570), .IN2(n4687), .IN3(g6782), .IN4(n2849), .Q(g30287) );
  AO22X1 U6043 ( .IN1(g1567), .IN2(n4317), .IN3(g1520), .IN4(n2849), .Q(g30279) );
  AO22X1 U6044 ( .IN1(g954), .IN2(n4693), .IN3(n2678), .IN4(g6368), .Q(g30670)
         );
  AO22X1 U6045 ( .IN1(g909), .IN2(n4693), .IN3(n4592), .IN4(n2746), .Q(g30638)
         );
  AO22X1 U6046 ( .IN1(g948), .IN2(n4692), .IN3(n2861), .IN4(n4591), .Q(g30271)
         );
  AO22X1 U6047 ( .IN1(test_so35), .IN2(n4323), .IN3(n2861), .IN4(n4592), .Q(
        g30265) );
  AO22X1 U6048 ( .IN1(g903), .IN2(n4692), .IN3(g6518), .IN4(n2907), .Q(g30249)
         );
  AO22X1 U6049 ( .IN1(g900), .IN2(n4323), .IN3(n4592), .IN4(n2907), .Q(g30247)
         );
  AO22X1 U6050 ( .IN1(g939), .IN2(n4692), .IN3(n2870), .IN4(g6518), .Q(g30264)
         );
  AO22X1 U6051 ( .IN1(g936), .IN2(n4693), .IN3(n2870), .IN4(g6368), .Q(g30259)
         );
  AO22X1 U6052 ( .IN1(g894), .IN2(n4692), .IN3(n4591), .IN4(n2845), .Q(g30293)
         );
  AO22X1 U6053 ( .IN1(g891), .IN2(n4693), .IN3(n4592), .IN4(n2845), .Q(g30286)
         );
  AO22X1 U6054 ( .IN1(g927), .IN2(n4693), .IN3(n2713), .IN4(n4592), .Q(g30649)
         );
  AO22X1 U6055 ( .IN1(g885), .IN2(n4692), .IN3(g6518), .IN4(n2665), .Q(g30681)
         );
  AO22X1 U6056 ( .IN1(g882), .IN2(n4693), .IN3(g6368), .IN4(n2665), .Q(g30676)
         );
  AO22X1 U6057 ( .IN1(g918), .IN2(n4693), .IN3(n2731), .IN4(n4592), .Q(g30643)
         );
  AO22X1 U6058 ( .IN1(g876), .IN2(n4692), .IN3(n4591), .IN4(n2856), .Q(g30277)
         );
  AO22X1 U6059 ( .IN1(g873), .IN2(n4693), .IN3(g6368), .IN4(n2856), .Q(g30269)
         );
  AO22X1 U6060 ( .IN1(g261), .IN2(n4697), .IN3(n2872), .IN4(n4593), .Q(g30263)
         );
  AO22X1 U6061 ( .IN1(g258), .IN2(n4698), .IN3(n2872), .IN4(g6231), .Q(g30258)
         );
  AO22X1 U6062 ( .IN1(g216), .IN2(n4697), .IN3(g6313), .IN4(n2925), .Q(g30246)
         );
  AO22X1 U6063 ( .IN1(g213), .IN2(n4698), .IN3(g138), .IN4(n2925), .Q(g30245)
         );
  AO22X1 U6064 ( .IN1(g252), .IN2(n4697), .IN3(n2878), .IN4(g6313), .Q(g30257)
         );
  AO22X1 U6065 ( .IN1(g249), .IN2(n4698), .IN3(n2878), .IN4(g138), .Q(g30254)
         );
  AO22X1 U6066 ( .IN1(g207), .IN2(n4697), .IN3(n4593), .IN4(n2850), .Q(g30284)
         );
  AO22X1 U6067 ( .IN1(g204), .IN2(n4318), .IN3(g6231), .IN4(n2850), .Q(g30276)
         );
  AO22X1 U6068 ( .IN1(g240), .IN2(n4318), .IN3(n2732), .IN4(g6231), .Q(g30641)
         );
  AO22X1 U6069 ( .IN1(g198), .IN2(n4697), .IN3(g6313), .IN4(n2679), .Q(g30674)
         );
  AO22X1 U6070 ( .IN1(g195), .IN2(n4698), .IN3(g138), .IN4(n2679), .Q(g30668)
         );
  AO22X1 U6071 ( .IN1(g231), .IN2(n4318), .IN3(n2747), .IN4(g6231), .Q(g30637)
         );
  AO22X1 U6072 ( .IN1(test_so13), .IN2(n4697), .IN3(n4593), .IN4(n2864), .Q(
        g30267) );
  AO22X1 U6073 ( .IN1(g186), .IN2(n4318), .IN3(g138), .IN4(n2864), .Q(g30261)
         );
  AO22X1 U6074 ( .IN1(g2318), .IN2(n4682), .IN3(n2680), .IN4(n4587), .Q(g30673) );
  AO22X1 U6075 ( .IN1(g2309), .IN2(n4682), .IN3(n2694), .IN4(n4587), .Q(g30666) );
  AO22X1 U6076 ( .IN1(g1624), .IN2(n4686), .IN3(n2695), .IN4(g6782), .Q(g30664) );
  AO22X1 U6077 ( .IN1(g1615), .IN2(n4686), .IN3(n2712), .IN4(n4589), .Q(g30657) );
  AO22X1 U6078 ( .IN1(g930), .IN2(n4312), .IN3(n2713), .IN4(n4591), .Q(g30655)
         );
  AO22X1 U6079 ( .IN1(g921), .IN2(n4312), .IN3(n2731), .IN4(n4591), .Q(g30648)
         );
  AO22X1 U6080 ( .IN1(g243), .IN2(n4696), .IN3(n2732), .IN4(n4593), .Q(g30646)
         );
  AO22X1 U6081 ( .IN1(g234), .IN2(n4696), .IN3(n2747), .IN4(n4593), .Q(g30640)
         );
  AO22X1 U6082 ( .IN1(g957), .IN2(n4312), .IN3(n2678), .IN4(g6518), .Q(g30677)
         );
  AO22X1 U6083 ( .IN1(g912), .IN2(n4312), .IN3(n4591), .IN4(n2746), .Q(g30642)
         );
  AO22X1 U6084 ( .IN1(g2394), .IN2(n4664), .IN3(n2796), .IN4(n4608), .Q(g30341) );
  AO22X1 U6085 ( .IN1(g2391), .IN2(n4664), .IN3(n2592), .IN4(n4608), .Q(g30709) );
  AO22X1 U6086 ( .IN1(g2388), .IN2(n4664), .IN3(n2964), .IN4(n4608), .Q(g29621) );
  AO22X1 U6087 ( .IN1(g1700), .IN2(n4667), .IN3(n2797), .IN4(n4620), .Q(g30503) );
  AO22X1 U6088 ( .IN1(g1697), .IN2(n4667), .IN3(n2593), .IN4(n4620), .Q(g30706) );
  AO22X1 U6089 ( .IN1(g1694), .IN2(n4667), .IN3(n2965), .IN4(n4620), .Q(g29617) );
  AO22X1 U6090 ( .IN1(g1006), .IN2(n4672), .IN3(n2798), .IN4(g6712), .Q(g30485) );
  AO22X1 U6091 ( .IN1(g1003), .IN2(n4672), .IN3(n2594), .IN4(g6712), .Q(g30703) );
  AO22X1 U6092 ( .IN1(g1000), .IN2(n4672), .IN3(n2969), .IN4(g6712), .Q(g29612) );
  AO22X1 U6093 ( .IN1(g2395), .IN2(n4663), .IN3(n2796), .IN4(n4606), .Q(g30356) );
  AO22X1 U6094 ( .IN1(g2393), .IN2(n4665), .IN3(n2796), .IN4(n4610), .Q(g30505) );
  AO22X1 U6095 ( .IN1(g2392), .IN2(n4663), .IN3(n2592), .IN4(n4606), .Q(g30566) );
  AO22X1 U6096 ( .IN1(g2390), .IN2(n4665), .IN3(n2592), .IN4(n4610), .Q(g30707) );
  AO22X1 U6097 ( .IN1(g2389), .IN2(n4663), .IN3(n2964), .IN4(n4606), .Q(g29623) );
  AO22X1 U6098 ( .IN1(g2387), .IN2(n4665), .IN3(n2964), .IN4(n4610), .Q(g29618) );
  AO22X1 U6099 ( .IN1(g1701), .IN2(n4666), .IN3(n2797), .IN4(n4618), .Q(g30338) );
  AO22X1 U6100 ( .IN1(g1699), .IN2(n4668), .IN3(n2797), .IN4(n4622), .Q(g30487) );
  AO22X1 U6101 ( .IN1(g1698), .IN2(n4666), .IN3(n2593), .IN4(n4618), .Q(g30708) );
  AO22X1 U6102 ( .IN1(g1696), .IN2(n4668), .IN3(n2593), .IN4(n4622), .Q(g30704) );
  AO22X1 U6103 ( .IN1(g1695), .IN2(n4666), .IN3(n2965), .IN4(n4618), .Q(g29620) );
  AO22X1 U6104 ( .IN1(g1693), .IN2(n4668), .IN3(n2965), .IN4(n4622), .Q(g29613) );
  AO22X1 U6105 ( .IN1(test_so39), .IN2(n4670), .IN3(n2798), .IN4(n4630), .Q(
        g30500) );
  AO22X1 U6106 ( .IN1(g1005), .IN2(n4674), .IN3(n2798), .IN4(g5472), .Q(g30470) );
  AO22X1 U6107 ( .IN1(g1004), .IN2(n4670), .IN3(n2594), .IN4(n4630), .Q(g30705) );
  AO22X1 U6108 ( .IN1(g1002), .IN2(n4674), .IN3(n2594), .IN4(g5472), .Q(g30701) );
  AO22X1 U6109 ( .IN1(g1001), .IN2(n4670), .IN3(n2969), .IN4(n4630), .Q(g29616) );
  AO22X1 U6110 ( .IN1(g999), .IN2(n4674), .IN3(n2969), .IN4(g5472), .Q(g29609)
         );
  AO22X1 U6111 ( .IN1(g320), .IN2(n4675), .IN3(n2799), .IN4(n4640), .Q(g30482)
         );
  AO22X1 U6112 ( .IN1(g319), .IN2(n4677), .IN3(n2799), .IN4(n4641), .Q(g30468)
         );
  AO22X1 U6113 ( .IN1(g318), .IN2(n4678), .IN3(n2799), .IN4(n4643), .Q(g30455)
         );
  AO22X1 U6114 ( .IN1(g317), .IN2(n4675), .IN3(n2615), .IN4(n4640), .Q(g30702)
         );
  AO22X1 U6115 ( .IN1(test_so18), .IN2(n4677), .IN3(n2615), .IN4(n4641), .Q(
        g30700) );
  AO22X1 U6116 ( .IN1(g315), .IN2(n4678), .IN3(n2615), .IN4(n4643), .Q(g30699)
         );
  AO22X1 U6117 ( .IN1(g314), .IN2(n4675), .IN3(n2973), .IN4(n4640), .Q(g29611)
         );
  AO22X1 U6118 ( .IN1(g313), .IN2(n4677), .IN3(n2973), .IN4(n4641), .Q(g29608)
         );
  AO22X1 U6119 ( .IN1(g312), .IN2(n4678), .IN3(n2973), .IN4(n4643), .Q(g29606)
         );
  AO22X1 U6120 ( .IN1(g2339), .IN2(n4367), .IN3(n2846), .IN4(n4679), .Q(g30297) );
  AO22X1 U6121 ( .IN1(g1645), .IN2(n4368), .IN3(n2853), .IN4(n4684), .Q(g30288) );
  AO22X1 U6122 ( .IN1(g264), .IN2(n4369), .IN3(n2872), .IN4(n4694), .Q(g30268)
         );
  AO22X1 U6123 ( .IN1(g2285), .IN2(n4680), .IN3(g2241), .IN4(n2840), .Q(g30304) );
  AO22X1 U6124 ( .IN1(g1591), .IN2(n4685), .IN3(g1547), .IN4(n2841), .Q(g30302) );
  AO22X1 U6125 ( .IN1(g915), .IN2(n4362), .IN3(n4690), .IN4(n2746), .Q(g30647)
         );
  AO22X1 U6126 ( .IN1(g897), .IN2(n4691), .IN3(n4690), .IN4(n2845), .Q(g30298)
         );
  AO22X1 U6127 ( .IN1(g210), .IN2(n4695), .IN3(g165), .IN4(n2850), .Q(g30292)
         );
  AO22X1 U6128 ( .IN1(g2294), .IN2(n4367), .IN3(g2241), .IN4(n2880), .Q(g30260) );
  AO22X1 U6129 ( .IN1(g2276), .IN2(n4367), .IN3(g2241), .IN4(n2656), .Q(g30695) );
  AO22X1 U6130 ( .IN1(g2267), .IN2(n4367), .IN3(g2241), .IN4(n2844), .Q(g30300) );
  AO22X1 U6131 ( .IN1(g1600), .IN2(n4368), .IN3(g1547), .IN4(n2886), .Q(g30255) );
  AO22X1 U6132 ( .IN1(g1582), .IN2(n4368), .IN3(g1547), .IN4(n2658), .Q(g30692) );
  AO22X1 U6133 ( .IN1(g1573), .IN2(n4368), .IN3(g1547), .IN4(n2849), .Q(g30294) );
  AO22X1 U6134 ( .IN1(g906), .IN2(n4691), .IN3(n4690), .IN4(n2907), .Q(g30251)
         );
  AO22X1 U6135 ( .IN1(g888), .IN2(n4691), .IN3(n4690), .IN4(n2665), .Q(g30687)
         );
  AO22X1 U6136 ( .IN1(g879), .IN2(n4691), .IN3(n4690), .IN4(n2856), .Q(g30285)
         );
  AO22X1 U6137 ( .IN1(g219), .IN2(n4369), .IN3(g165), .IN4(n2925), .Q(g30248)
         );
  AO22X1 U6138 ( .IN1(g201), .IN2(n4369), .IN3(g165), .IN4(n2679), .Q(g30680)
         );
  AO22X1 U6139 ( .IN1(g192), .IN2(n4369), .IN3(g165), .IN4(n2864), .Q(g30275)
         );
  ISOLANDX1 U6140 ( .D(g3002), .ISO(n4066), .Q(n4065) );
  INVX0 U6141 ( .IN(g2214), .QN(n4683) );
  INVX0 U6142 ( .IN(g6368), .QN(n4693) );
  INVX0 U6143 ( .IN(g7084), .QN(n4681) );
  INVX0 U6144 ( .IN(g6782), .QN(n4687) );
  INVX0 U6145 ( .IN(g6518), .QN(n4692) );
  INVX0 U6146 ( .IN(g6313), .QN(n4697) );
  INVX0 U6147 ( .IN(g1520), .QN(n4688) );
  INVX0 U6148 ( .IN(g138), .QN(n4698) );
  OAI222X1 U6149 ( .IN1(n4324), .IN2(g2209), .IN3(n4367), .IN4(g2208), .IN5(
        n4681), .IN6(g2210), .QN(n3877) );
  OAI222X1 U6150 ( .IN1(n4324), .IN2(g2206), .IN3(n4367), .IN4(g2205), .IN5(
        n4681), .IN6(g2207), .QN(n3878) );
  OAI222X1 U6151 ( .IN1(n4324), .IN2(g2218), .IN3(n4682), .IN4(g2219), .IN5(
        n4367), .IN6(g2217), .QN(n3879) );
  OAI222X1 U6152 ( .IN1(n4688), .IN2(test_so52), .IN3(n4368), .IN4(g1514), 
        .IN5(n4687), .IN6(g1516), .QN(n3774) );
  OAI222X1 U6153 ( .IN1(n4317), .IN2(g1512), .IN3(n4368), .IN4(g1511), .IN5(
        n4687), .IN6(g1513), .QN(n3775) );
  OAI222X1 U6154 ( .IN1(n4317), .IN2(g1524), .IN3(n4687), .IN4(g1525), .IN5(
        n4368), .IN6(g1523), .QN(n3776) );
  OAI222X1 U6155 ( .IN1(n4323), .IN2(g821), .IN3(n4691), .IN4(g820), .IN5(
        n4692), .IN6(g822), .QN(n3804) );
  OAI222X1 U6156 ( .IN1(n4323), .IN2(g818), .IN3(n4691), .IN4(g817), .IN5(
        n4692), .IN6(g819), .QN(n3805) );
  OAI222X1 U6157 ( .IN1(n4323), .IN2(g830), .IN3(n4692), .IN4(g831), .IN5(
        n4691), .IN6(g829), .QN(n3806) );
  OAI222X1 U6158 ( .IN1(n4698), .IN2(g133), .IN3(n4369), .IN4(g132), .IN5(
        n4697), .IN6(g134), .QN(n3832) );
  OAI222X1 U6159 ( .IN1(n4318), .IN2(g130), .IN3(n4369), .IN4(g129), .IN5(
        n4697), .IN6(g131), .QN(n3833) );
  OAI222X1 U6160 ( .IN1(n4318), .IN2(g142), .IN3(n4697), .IN4(g143), .IN5(
        n4369), .IN6(g141), .QN(n3834) );
  OAI222X1 U6161 ( .IN1(n4324), .IN2(g2233), .IN3(n4681), .IN4(g2234), .IN5(
        n4367), .IN6(g2232), .QN(n3872) );
  OAI222X1 U6162 ( .IN1(n4324), .IN2(g2224), .IN3(n4681), .IN4(test_so74), 
        .IN5(n4367), .IN6(g2223), .QN(n3871) );
  OAI222X1 U6163 ( .IN1(n4324), .IN2(g2221), .IN3(n4682), .IN4(g2222), .IN5(
        n4367), .IN6(g2220), .QN(n3873) );
  OAI222X1 U6164 ( .IN1(n4688), .IN2(g1539), .IN3(n4687), .IN4(g1540), .IN5(
        n4368), .IN6(g1538), .QN(n3769) );
  OAI222X1 U6165 ( .IN1(n4688), .IN2(g1530), .IN3(n4687), .IN4(g1531), .IN5(
        n4368), .IN6(g1529), .QN(n3768) );
  OAI222X1 U6166 ( .IN1(n4688), .IN2(g1527), .IN3(n4687), .IN4(g1528), .IN5(
        n4368), .IN6(g1526), .QN(n3770) );
  OAI222X1 U6167 ( .IN1(n4323), .IN2(g845), .IN3(n4692), .IN4(g846), .IN5(
        n4691), .IN6(g844), .QN(n3799) );
  OAI222X1 U6168 ( .IN1(n4323), .IN2(g836), .IN3(n4692), .IN4(g837), .IN5(
        n4691), .IN6(g835), .QN(n3798) );
  OAI222X1 U6169 ( .IN1(n4693), .IN2(g833), .IN3(n4692), .IN4(g834), .IN5(
        n4691), .IN6(g832), .QN(n3800) );
  OAI222X1 U6170 ( .IN1(n4698), .IN2(g157), .IN3(n4697), .IN4(g158), .IN5(
        n4369), .IN6(g156), .QN(n3827) );
  OAI222X1 U6171 ( .IN1(n4698), .IN2(g148), .IN3(n4697), .IN4(g149), .IN5(
        n4369), .IN6(g147), .QN(n3826) );
  OAI222X1 U6172 ( .IN1(n4698), .IN2(g145), .IN3(n4697), .IN4(g146), .IN5(
        n4369), .IN6(test_so11), .QN(n3828) );
  OA22X1_S38584 U6173 ( .IN1(g2451), .IN2(n1619), .IN3(n3524), .IN4(n3513), .Q(g27334) );
  OA22X1_S38584 U6174 ( .IN1(g2448), .IN2(n1618), .IN3(n3524), .IN4(n3523), .Q(g27323) );
  OA22X1_S38584 U6175 ( .IN1(g2459), .IN2(n1617), .IN3(n3524), .IN4(n3538), .Q(g27309) );
  OA22X1_S38584 U6176 ( .IN1(g1757), .IN2(n1616), .IN3(n3550), .IN4(n3530), .Q(g27317) );
  OA22X1_S38584 U6177 ( .IN1(g1754), .IN2(n1615), .IN3(n3550), .IN4(n3549), .Q(g27303) );
  OA22X1_S38584 U6178 ( .IN1(g1765), .IN2(n1614), .IN3(n3550), .IN4(n3573), .Q(g27289) );
  OA22X1_S38584 U6179 ( .IN1(g1063), .IN2(n1613), .IN3(n3585), .IN4(n3556), .Q(g27297) );
  OA22X1_S38584 U6180 ( .IN1(g1060), .IN2(n1612), .IN3(n3585), .IN4(n3584), .Q(g27283) );
  OA22X1_S38584 U6181 ( .IN1(test_so37), .IN2(n1611), .IN3(n3585), .IN4(n3609), .Q(
        g27272) );
  OA22X1_S38584 U6182 ( .IN1(g376), .IN2(n1610), .IN3(n3621), .IN4(n3591), .Q(g27277)
         );
  OA22X1_S38584 U6183 ( .IN1(g373), .IN2(n1609), .IN3(n3621), .IN4(n3620), .Q(g27266)
         );
  OA22X1_S38584 U6184 ( .IN1(g384), .IN2(n1608), .IN3(n3621), .IN4(n3643), .Q(g27260)
         );
  OA22X1_S38584 U6185 ( .IN1(g2398), .IN2(n3031), .IN3(n4664), .IN4(n3029), .Q(g29185) );
  NOR2X0 U6186 ( .IN1(n3030), .IN2(n4524), .QN(n3031) );
  OA22X1_S38584 U6187 ( .IN1(g1704), .IN2(n3063), .IN3(n4667), .IN4(n3033), .Q(g29181) );
  NOR2X0 U6188 ( .IN1(n3034), .IN2(n4525), .QN(n3063) );
  OA22X1_S38584 U6189 ( .IN1(g1010), .IN2(n3095), .IN3(n4672), .IN4(n3065), .Q(g29173) );
  NOR2X0 U6190 ( .IN1(n3066), .IN2(n4671), .QN(n3095) );
  OA22X1_S38584 U6191 ( .IN1(g2396), .IN2(n3028), .IN3(n4663), .IN4(n3029), .Q(g29187) );
  NOR2X0 U6192 ( .IN1(n3030), .IN2(n4509), .QN(n3028) );
  OA22X1_S38584 U6193 ( .IN1(g2397), .IN2(n3035), .IN3(n4665), .IN4(n3029), .Q(g29182) );
  NOR2X0 U6194 ( .IN1(n3030), .IN2(n4516), .QN(n3035) );
  OA22X1_S38584 U6195 ( .IN1(g1702), .IN2(n3032), .IN3(n4666), .IN4(n3033), .Q(g29184) );
  NOR2X0 U6196 ( .IN1(n3034), .IN2(n4511), .QN(n3032) );
  OA22X1_S38584 U6197 ( .IN1(g1703), .IN2(n3067), .IN3(n4668), .IN4(n3033), .Q(g29178) );
  NOR2X0 U6198 ( .IN1(n3034), .IN2(n4518), .QN(n3067) );
  OA22X1_S38584 U6199 ( .IN1(g1008), .IN2(n3064), .IN3(n4670), .IN4(n3065), .Q(g29179) );
  NOR2X0 U6200 ( .IN1(n3066), .IN2(n4669), .QN(n3064) );
  OA22X1_S38584 U6201 ( .IN1(g1009), .IN2(n3099), .IN3(n4674), .IN4(n3065), .Q(g29170) );
  NOR2X0 U6202 ( .IN1(n3066), .IN2(n4673), .QN(n3099) );
  OA22X1_S38584 U6203 ( .IN1(g321), .IN2(n3096), .IN3(n4675), .IN4(n3097), .Q(g29172)
         );
  NOR2X0 U6204 ( .IN1(n3098), .IN2(n4506), .QN(n3096) );
  OA22X1_S38584 U6205 ( .IN1(g323), .IN2(n3126), .IN3(n4677), .IN4(n3097), .Q(g29169)
         );
  NOR2X0 U6206 ( .IN1(n3098), .IN2(n4676), .QN(n3126) );
  OA22X1_S38584 U6207 ( .IN1(g322), .IN2(n3127), .IN3(n4678), .IN4(n3097), .Q(g29167)
         );
  NOR2X0 U6208 ( .IN1(n3098), .IN2(n4520), .QN(n3127) );
  INVX0 U6209 ( .IN(g6782), .QN(n4686) );
  INVX0 U6210 ( .IN(g6313), .QN(n4696) );
  NBUFFX2 U6211 ( .IN(g2625), .Q(g7390) );
  NBUFFX2 U6212 ( .IN(g1931), .Q(g7194) );
  NBUFFX2 U6213 ( .IN(g1237), .Q(g6944) );
  NBUFFX2 U6214 ( .IN(g551), .Q(g6642) );
  NOR4X0 U6215 ( .IN1(n3867), .IN2(n3868), .IN3(n3869), .IN4(n3870), .QN(n3866) );
  XOR2X1 U6216 ( .IN1(n3873), .IN2(g2180), .Q(n3868) );
  XOR2X1 U6217 ( .IN1(n3871), .IN2(g2185), .Q(n3870) );
  XOR2X1 U6218 ( .IN1(n3872), .IN2(g2200), .Q(n3869) );
  NOR4X0 U6219 ( .IN1(n3764), .IN2(n3765), .IN3(n3766), .IN4(n3767), .QN(n3763) );
  XOR2X1 U6220 ( .IN1(n3770), .IN2(g1486), .Q(n3765) );
  XOR2X1 U6221 ( .IN1(n3768), .IN2(g1491), .Q(n3767) );
  XOR2X1 U6222 ( .IN1(n3769), .IN2(g1506), .Q(n3766) );
  NOR4X0 U6223 ( .IN1(n3794), .IN2(n3795), .IN3(n3796), .IN4(n3797), .QN(n3793) );
  XOR2X1 U6224 ( .IN1(n3800), .IN2(g797), .Q(n3795) );
  XOR2X1 U6225 ( .IN1(n3798), .IN2(g801), .Q(n3797) );
  XOR2X1 U6226 ( .IN1(n3799), .IN2(g813), .Q(n3796) );
  NOR4X0 U6227 ( .IN1(n3822), .IN2(n3823), .IN3(n3824), .IN4(n3825), .QN(n3821) );
  XOR2X1 U6228 ( .IN1(n3828), .IN2(g109), .Q(n3823) );
  XOR2X1 U6229 ( .IN1(n3826), .IN2(g113), .Q(n3825) );
  XOR2X1 U6230 ( .IN1(n3827), .IN2(g125), .Q(n3824) );
  NBUFFX2 U6231 ( .IN(g2619), .Q(n4604) );
  XOR2X1 U6232 ( .IN1(n4554), .IN2(n4555), .Q(n3881) );
  OA222X1 U6233 ( .IN1(n4324), .IN2(g2227), .IN3(n4682), .IN4(g2228), .IN5(
        n4367), .IN6(g2226), .Q(n4554) );
  XOR2X1 U6234 ( .IN1(n4556), .IN2(n4557), .Q(n3778) );
  OA222X1 U6235 ( .IN1(n4317), .IN2(g1533), .IN3(n4687), .IN4(g1534), .IN5(
        n4368), .IN6(g1532), .Q(n4556) );
  XOR2X1 U6236 ( .IN1(n4558), .IN2(n4559), .Q(n3808) );
  OA222X1 U6237 ( .IN1(n4323), .IN2(test_so32), .IN3(n4692), .IN4(g840), .IN5(
        n4691), .IN6(g838), .Q(n4558) );
  XOR2X1 U6238 ( .IN1(n4560), .IN2(n4561), .Q(n3836) );
  OA222X1 U6239 ( .IN1(n4318), .IN2(g151), .IN3(n4697), .IN4(g152), .IN5(n4369), .IN6(g150), .Q(n4560) );
  XOR2X1 U6240 ( .IN1(n4562), .IN2(n4563), .Q(n3880) );
  OA222X1 U6241 ( .IN1(n4324), .IN2(g2230), .IN3(n4682), .IN4(g2231), .IN5(
        n4367), .IN6(g2229), .Q(n4562) );
  XOR2X1 U6242 ( .IN1(n4564), .IN2(n4565), .Q(n3777) );
  OA222X1 U6243 ( .IN1(n4688), .IN2(g1536), .IN3(n4687), .IN4(test_so53), 
        .IN5(n4368), .IN6(g1535), .Q(n4564) );
  XOR2X1 U6244 ( .IN1(n4566), .IN2(n4567), .Q(n3807) );
  OA222X1 U6245 ( .IN1(n4323), .IN2(g842), .IN3(n4692), .IN4(g843), .IN5(n4691), .IN6(g841), .Q(n4566) );
  XOR2X1 U6246 ( .IN1(n4568), .IN2(n4569), .Q(n3835) );
  OA222X1 U6247 ( .IN1(n4698), .IN2(g154), .IN3(n4697), .IN4(g155), .IN5(n4369), .IN6(g153), .Q(n4568) );
  NBUFFX2 U6248 ( .IN(g2624), .Q(n4599) );
  NBUFFX2 U6249 ( .IN(g1930), .Q(n4611) );
  NBUFFX2 U6250 ( .IN(g1236), .Q(n4623) );
  NBUFFX2 U6251 ( .IN(g550), .Q(n4633) );
  NBUFFX2 U6252 ( .IN(g3080), .Q(n4597) );
  INVX0 U6253 ( .IN(g7084), .QN(n4682) );
  NBUFFX2 U6254 ( .IN(g1088), .Q(n4629) );
  NOR2X0 U6255 ( .IN1(n1606), .IN2(n2992), .QN(g29357) );
  XOR2X1 U6256 ( .IN1(n2982), .IN2(g2124), .Q(n2992) );
  NOR2X0 U6257 ( .IN1(n1605), .IN2(n2993), .QN(g29355) );
  XOR2X1 U6258 ( .IN1(n2985), .IN2(g1430), .Q(n2993) );
  NOR2X0 U6259 ( .IN1(n1604), .IN2(n2994), .QN(g29354) );
  XOR2X1 U6260 ( .IN1(n2988), .IN2(g744), .Q(n2994) );
  NOR2X0 U6261 ( .IN1(n1603), .IN2(n2995), .QN(g29353) );
  XOR2X1 U6262 ( .IN1(n2991), .IN2(g56), .Q(n2995) );
  NAND4X0 U6263 ( .IN1(n3898), .IN2(n3899), .IN3(n3900), .IN4(n3901), .QN(
        g26149) );
  OA221X1 U6264 ( .IN1(n3902), .IN2(n4441), .IN3(n3903), .IN4(n4338), .IN5(
        n3904), .Q(n3901) );
  OA221X1 U6265 ( .IN1(n3916), .IN2(DFF_149_n1), .IN3(n3917), .IN4(n4436), 
        .IN5(n3918), .Q(n3898) );
  OA221X1 U6266 ( .IN1(n3912), .IN2(n4444), .IN3(n3913), .IN4(n4339), .IN5(
        n3914), .Q(n3899) );
  AND4X1 U6267 ( .IN1(n1607), .IN2(g2883), .IN3(g2924), .IN4(n4222), .Q(g13110) );
  NOR4X0 U6268 ( .IN1(g2920), .IN2(g2917), .IN3(g2912), .IN4(g2888), .QN(n4222) );
  AO221X1 U6269 ( .IN1(g3110), .IN2(n1746), .IN3(n1745), .IN4(DFF_144_n1), 
        .IN5(n1574), .Q(g25435) );
  AO21X1 U6270 ( .IN1(n1745), .IN2(DFF_146_n1), .IN3(n1574), .Q(g24734) );
  OA222X1 U6271 ( .IN1(n4370), .IN2(g2651), .IN3(n4299), .IN4(g2649), .IN5(
        n4314), .IN6(g2650), .Q(n3275) );
  OA222X1 U6272 ( .IN1(n4315), .IN2(g1957), .IN3(n4366), .IN4(g1955), .IN5(
        n4296), .IN6(g1956), .Q(n3316) );
  OA222X1 U6273 ( .IN1(n4316), .IN2(g1263), .IN3(n4300), .IN4(g1261), .IN5(
        n4371), .IN6(g1262), .Q(n3356) );
  OA222X1 U6274 ( .IN1(n4372), .IN2(g577), .IN3(n4313), .IN4(g575), .IN5(n4298), .IN6(g576), .Q(n3395) );
  INVX0 U6275 ( .IN(n4585), .QN(n4586) );
  INVX0 U6276 ( .IN(g51), .QN(n4585) );
  AO222X1 U6277 ( .IN1(g2495), .IN2(n4608), .IN3(g2498), .IN4(n4606), .IN5(
        g2492), .IN6(n4610), .Q(n4285) );
  AO222X1 U6278 ( .IN1(g1801), .IN2(n4620), .IN3(g1804), .IN4(n4618), .IN5(
        g1798), .IN6(n4622), .Q(n4284) );
  AO222X1 U6279 ( .IN1(g1104), .IN2(g5472), .IN3(g1110), .IN4(n4630), .IN5(
        g1107), .IN6(g6712), .Q(n4283) );
  AO222X1 U6280 ( .IN1(g420), .IN2(n4641), .IN3(g423), .IN4(n4640), .IN5(g417), 
        .IN6(n4643), .Q(n4282) );
  AO222X1 U6281 ( .IN1(g2456), .IN2(g5796), .IN3(g2458), .IN4(g2412), .IN5(
        g2454), .IN6(g5747), .Q(n3276) );
  AO222X1 U6282 ( .IN1(g1762), .IN2(g5738), .IN3(g1764), .IN4(g1718), .IN5(
        g1760), .IN6(g5695), .Q(n3317) );
  AO222X1 U6283 ( .IN1(g1068), .IN2(g5686), .IN3(g1070), .IN4(g1024), .IN5(
        g1066), .IN6(g5657), .Q(n3357) );
  AO222X1 U6284 ( .IN1(g381), .IN2(g5648), .IN3(g383), .IN4(g337), .IN5(g379), 
        .IN6(g5629), .Q(n3396) );
  OA222X1 U6285 ( .IN1(n4370), .IN2(g2654), .IN3(n4299), .IN4(g2652), .IN5(
        n4314), .IN6(g2653), .Q(n3288) );
  OA222X1 U6286 ( .IN1(n4315), .IN2(g1960), .IN3(n4366), .IN4(g1958), .IN5(
        n4296), .IN6(g1959), .Q(n3329) );
  OA222X1 U6287 ( .IN1(n4316), .IN2(g1266), .IN3(n4300), .IN4(g1264), .IN5(
        n4371), .IN6(g1265), .Q(n3369) );
  OA222X1 U6288 ( .IN1(n4372), .IN2(test_so25), .IN3(n4313), .IN4(g578), .IN5(
        n4298), .IN6(g579), .Q(n3408) );
  AO221X1 U6289 ( .IN1(g3112), .IN2(n1746), .IN3(test_so9), .IN4(n1745), .IN5(
        n1574), .Q(g25420) );
  AO221X1 U6290 ( .IN1(g3111), .IN2(n1746), .IN3(g3124), .IN4(n1745), .IN5(
        n1574), .Q(g25442) );
  AO222X1 U6291 ( .IN1(g2516), .IN2(n4608), .IN3(g2519), .IN4(n4606), .IN5(
        g2513), .IN6(n4610), .Q(n3448) );
  AO222X1 U6292 ( .IN1(g1822), .IN2(n4620), .IN3(test_so59), .IN4(n4618), 
        .IN5(g1819), .IN6(n4622), .Q(n3460) );
  AO222X1 U6293 ( .IN1(g1125), .IN2(g5472), .IN3(g1131), .IN4(n4630), .IN5(
        g1128), .IN6(g6712), .Q(n3472) );
  AO222X1 U6294 ( .IN1(g441), .IN2(n4641), .IN3(g444), .IN4(n4640), .IN5(g438), 
        .IN6(n4643), .Q(n3481) );
  NAND2X0 U6295 ( .IN1(g2257), .IN2(n4679), .QN(n4169) );
  NAND2X0 U6296 ( .IN1(g1563), .IN2(n4684), .QN(n4171) );
  NAND2X0 U6297 ( .IN1(g869), .IN2(n4689), .QN(n4174) );
  NAND2X0 U6298 ( .IN1(g181), .IN2(n4694), .QN(n4177) );
  OA222X1 U6299 ( .IN1(n4524), .IN2(g2418), .IN3(n4509), .IN4(g2421), .IN5(
        n4516), .IN6(g2429), .Q(n3542) );
  OA222X1 U6300 ( .IN1(n4525), .IN2(g1724), .IN3(n4511), .IN4(g1727), .IN5(
        n4518), .IN6(g1735), .Q(n3577) );
  OA222X1 U6301 ( .IN1(n4673), .IN2(g1041), .IN3(n4669), .IN4(g1033), .IN5(
        n4671), .IN6(g1030), .Q(n3613) );
  OA222X1 U6302 ( .IN1(n4676), .IN2(g343), .IN3(n4506), .IN4(test_so16), .IN5(
        n4520), .IN6(g354), .Q(n3647) );
  OA222X1 U6303 ( .IN1(n4370), .IN2(g2660), .IN3(n4299), .IN4(g2658), .IN5(
        n4314), .IN6(g2659), .Q(n3273) );
  OA222X1 U6304 ( .IN1(n4315), .IN2(g1966), .IN3(n4366), .IN4(g1964), .IN5(
        n4296), .IN6(test_so67), .Q(n3314) );
  OA222X1 U6305 ( .IN1(n4316), .IN2(g1272), .IN3(n4300), .IN4(g1270), .IN5(
        n4371), .IN6(g1271), .Q(n3354) );
  OA222X1 U6306 ( .IN1(n4372), .IN2(g586), .IN3(n4313), .IN4(g584), .IN5(n4298), .IN6(g585), .Q(n3393) );
  AO222X1 U6307 ( .IN1(g2426), .IN2(g5796), .IN3(g2428), .IN4(g2412), .IN5(
        g2424), .IN6(g5747), .Q(n3265) );
  AO222X1 U6308 ( .IN1(g1732), .IN2(g5738), .IN3(g1734), .IN4(g1718), .IN5(
        g1730), .IN6(g5695), .Q(n3306) );
  AO222X1 U6309 ( .IN1(g1038), .IN2(g5686), .IN3(g1040), .IN4(g1024), .IN5(
        g1036), .IN6(g5657), .Q(n3346) );
  AO222X1 U6310 ( .IN1(g351), .IN2(g5648), .IN3(g353), .IN4(g337), .IN5(g349), 
        .IN6(g5629), .Q(n3385) );
  AO222X1 U6311 ( .IN1(g2568), .IN2(n4602), .IN3(g2571), .IN4(n4600), .IN5(
        g2565), .IN6(n4604), .Q(n3843) );
  AO222X1 U6312 ( .IN1(g1874), .IN2(n4614), .IN3(g1877), .IN4(n4612), .IN5(
        test_so68), .IN6(n4616), .Q(n3845) );
  AO222X1 U6313 ( .IN1(g1180), .IN2(n4626), .IN3(g1183), .IN4(n4624), .IN5(
        test_so47), .IN6(n4628), .Q(n3847) );
  AO222X1 U6314 ( .IN1(g493), .IN2(n4636), .IN3(g496), .IN4(n4634), .IN5(g490), 
        .IN6(g6485), .Q(n3848) );
  AO222X1 U6315 ( .IN1(g1777), .IN2(g5738), .IN3(g1705), .IN4(g1718), .IN5(
        g1775), .IN6(g5695), .Q(n3311) );
  AO222X1 U6316 ( .IN1(g1083), .IN2(g5686), .IN3(g1011), .IN4(g1024), .IN5(
        g1081), .IN6(g5657), .Q(n3351) );
  AO222X1 U6317 ( .IN1(g396), .IN2(g5648), .IN3(g324), .IN4(g337), .IN5(g394), 
        .IN6(g5629), .Q(n3390) );
  AO222X1 U6318 ( .IN1(g2507), .IN2(n4608), .IN3(g2510), .IN4(n4606), .IN5(
        g2504), .IN6(n4610), .Q(n3447) );
  AO222X1 U6319 ( .IN1(g1813), .IN2(n4620), .IN3(g1816), .IN4(n4618), .IN5(
        g1810), .IN6(n4622), .Q(n3459) );
  AO222X1 U6320 ( .IN1(g432), .IN2(n4641), .IN3(g435), .IN4(n4640), .IN5(g429), 
        .IN6(n4643), .Q(n3480) );
  AO222X1 U6321 ( .IN1(g1116), .IN2(g5472), .IN3(g1122), .IN4(n4630), .IN5(
        test_so38), .IN6(g6712), .Q(n3471) );
  OA222X1 U6322 ( .IN1(n4664), .IN2(g2448), .IN3(n4509), .IN4(g2451), .IN5(
        n4516), .IN6(g2459), .Q(n3625) );
  OA222X1 U6323 ( .IN1(n4667), .IN2(g1754), .IN3(n4511), .IN4(g1757), .IN5(
        n4518), .IN6(g1765), .Q(n3652) );
  OA222X1 U6324 ( .IN1(n4673), .IN2(test_so37), .IN3(n4669), .IN4(g1063), 
        .IN5(n4671), .IN6(g1060), .Q(n3670) );
  OA222X1 U6325 ( .IN1(n4676), .IN2(g373), .IN3(n4506), .IN4(g376), .IN5(n4520), .IN6(g384), .Q(n3677) );
  OA222X1 U6326 ( .IN1(n4524), .IN2(g2433), .IN3(n4509), .IN4(g2436), .IN5(
        n4516), .IN6(g2444), .Q(n3567) );
  OA222X1 U6327 ( .IN1(n4525), .IN2(g1739), .IN3(n4511), .IN4(g1742), .IN5(
        n4518), .IN6(g1750), .Q(n3603) );
  OA222X1 U6328 ( .IN1(n4673), .IN2(g1056), .IN3(n4669), .IN4(g1048), .IN5(
        n4672), .IN6(g1045), .Q(n3637) );
  OA222X1 U6329 ( .IN1(n4676), .IN2(g358), .IN3(n4506), .IN4(g361), .IN5(n4520), .IN6(g369), .Q(n3664) );
  OA222X1 U6330 ( .IN1(n4524), .IN2(g2463), .IN3(n4509), .IN4(g2466), .IN5(
        n4516), .IN6(g2473), .Q(n3566) );
  OA222X1 U6331 ( .IN1(n4525), .IN2(test_so58), .IN3(n4511), .IN4(g1772), 
        .IN5(n4518), .IN6(g1779), .Q(n3602) );
  OA222X1 U6332 ( .IN1(n4673), .IN2(g1085), .IN3(n4669), .IN4(g1078), .IN5(
        n4671), .IN6(g1075), .Q(n3636) );
  OA222X1 U6333 ( .IN1(n4676), .IN2(g388), .IN3(n4506), .IN4(g391), .IN5(n4520), .IN6(g398), .Q(n3663) );
  OA222X1 U6334 ( .IN1(n4664), .IN2(g2503), .IN3(n4663), .IN4(g2501), .IN5(
        n4665), .IN6(g2502), .Q(n3004) );
  OA222X1 U6335 ( .IN1(n4667), .IN2(g1809), .IN3(n4666), .IN4(g1807), .IN5(
        n4668), .IN6(g1808), .Q(n3012) );
  OA222X1 U6336 ( .IN1(n4674), .IN2(g1114), .IN3(n4670), .IN4(g1113), .IN5(
        n4672), .IN6(g1115), .Q(n3020) );
  OA222X1 U6337 ( .IN1(n4677), .IN2(g428), .IN3(n4675), .IN4(g426), .IN5(n4678), .IN6(test_so17), .Q(n3027) );
  AO21X1 U6338 ( .IN1(g5388), .IN2(DFF_1612_n1), .IN3(n4365), .Q(g16496) );
  OA222X1 U6339 ( .IN1(n4524), .IN2(g2524), .IN3(n4509), .IN4(test_so81), 
        .IN5(n4516), .IN6(g2523), .Q(n3444) );
  OA222X1 U6340 ( .IN1(n4525), .IN2(g1830), .IN3(n4511), .IN4(g1828), .IN5(
        n4518), .IN6(g1829), .Q(n3456) );
  OA222X1 U6341 ( .IN1(n4673), .IN2(g1135), .IN3(n4669), .IN4(g1134), .IN5(
        n4671), .IN6(g1136), .Q(n3468) );
  OA222X1 U6342 ( .IN1(n4676), .IN2(g449), .IN3(n4506), .IN4(g447), .IN5(n4520), .IN6(g448), .Q(n3477) );
  AO221X1 U6343 ( .IN1(n4077), .IN2(test_so88), .IN3(g2670), .IN4(n4604), 
        .IN5(n4078), .Q(n3256) );
  AO22X1 U6344 ( .IN1(g2673), .IN2(n4602), .IN3(g2676), .IN4(n4600), .Q(n4078)
         );
  NOR2X0 U6345 ( .IN1(g12499), .IN2(n4384), .QN(n4077) );
  AO221X1 U6346 ( .IN1(n4083), .IN2(g1922), .IN3(g1976), .IN4(n4616), .IN5(
        n4084), .Q(n3297) );
  AO22X1 U6347 ( .IN1(g1979), .IN2(n4614), .IN3(g1982), .IN4(n4612), .Q(n4084)
         );
  NOR2X0 U6348 ( .IN1(g12482), .IN2(n4384), .QN(n4083) );
  AO221X1 U6349 ( .IN1(n4089), .IN2(test_so45), .IN3(g1282), .IN4(n4628), 
        .IN5(n4090), .Q(n3338) );
  AO22X1 U6350 ( .IN1(g1285), .IN2(n4626), .IN3(g1288), .IN4(n4624), .Q(n4090)
         );
  NOR2X0 U6351 ( .IN1(g12467), .IN2(n4384), .QN(n4089) );
  AO221X1 U6352 ( .IN1(n4094), .IN2(g542), .IN3(g596), .IN4(g6485), .IN5(n4095), .Q(n3378) );
  AO22X1 U6353 ( .IN1(g599), .IN2(n4636), .IN3(g602), .IN4(n4634), .Q(n4095)
         );
  NOR2X0 U6354 ( .IN1(g12457), .IN2(n4384), .QN(n4094) );
  AO221X1 U6355 ( .IN1(g2661), .IN2(g7302), .IN3(n4081), .IN4(g2598), .IN5(
        n4082), .Q(n3257) );
  AO22X1 U6356 ( .IN1(g2664), .IN2(n4602), .IN3(g2667), .IN4(n4600), .Q(n4082)
         );
  NOR2X0 U6357 ( .IN1(g12539), .IN2(n4384), .QN(n4081) );
  AO221X1 U6358 ( .IN1(g1967), .IN2(g7052), .IN3(n4087), .IN4(g1904), .IN5(
        n4088), .Q(n3298) );
  AO22X1 U6359 ( .IN1(g1970), .IN2(n4614), .IN3(g1973), .IN4(n4612), .Q(n4088)
         );
  NOR2X0 U6360 ( .IN1(g12524), .IN2(n4384), .QN(n4087) );
  AO221X1 U6361 ( .IN1(g1273), .IN2(g6750), .IN3(n4092), .IN4(g1210), .IN5(
        n4093), .Q(n3339) );
  AO22X1 U6362 ( .IN1(g1276), .IN2(n4626), .IN3(g1279), .IN4(n4624), .Q(n4093)
         );
  NOR2X0 U6363 ( .IN1(g12507), .IN2(n4384), .QN(n4092) );
  AO221X1 U6364 ( .IN1(g587), .IN2(n4638), .IN3(n4096), .IN4(g524), .IN5(n4097), .Q(n3379) );
  AO22X1 U6365 ( .IN1(g590), .IN2(n4636), .IN3(g593), .IN4(n4634), .Q(n4097)
         );
  NOR2X0 U6366 ( .IN1(g12487), .IN2(n4384), .QN(n4096) );
  AO21X1 U6367 ( .IN1(n4125), .IN2(n1587), .IN3(n1586), .Q(n2481) );
  NAND4X0 U6368 ( .IN1(g2920), .IN2(g2912), .IN3(n4479), .IN4(n4349), .QN(
        n4125) );
  OAI22X1 U6369 ( .IN1(n4570), .IN2(n4571), .IN3(n4572), .IN4(g506), .QN(n3855) );
  OR2X1 U6370 ( .IN1(n4636), .IN2(g16297), .Q(n4572) );
  XOR2X1 U6371 ( .IN1(n4202), .IN2(n4203), .Q(n4201) );
  XOR3X1 U6372 ( .IN1(g2975), .IN2(g2972), .IN3(n4204), .Q(n4203) );
  XNOR3X1 U6373 ( .IN1(n4205), .IN2(g2963), .IN3(g2874), .Q(n4202) );
  XOR2X1 U6374 ( .IN1(g2981), .IN2(g2978), .Q(n4204) );
  XOR2X1 U6375 ( .IN1(n4213), .IN2(n4214), .Q(n4212) );
  XOR3X1 U6376 ( .IN1(g2953), .IN2(g2947), .IN3(n4215), .Q(n4214) );
  XNOR3X1 U6377 ( .IN1(n4216), .IN2(g2938), .IN3(g2935), .Q(n4213) );
  XOR2X1 U6378 ( .IN1(g2959), .IN2(g2956), .Q(n4215) );
  AO21X1 U6379 ( .IN1(g1192), .IN2(DFF_783_n1), .IN3(n3854), .Q(n3174) );
  OA221X1 U6380 ( .IN1(n4626), .IN2(DFF_792_n1), .IN3(n4316), .IN4(n3855), 
        .IN5(n4454), .Q(n3854) );
  NAND2X0 U6381 ( .IN1(test_so79), .IN2(n3192), .QN(n3003) );
  NAND2X0 U6382 ( .IN1(g1690), .IN2(n3208), .QN(n3011) );
  NAND2X0 U6383 ( .IN1(g996), .IN2(n3221), .QN(n3019) );
  NAND2X0 U6384 ( .IN1(g309), .IN2(n3233), .QN(n3026) );
  NAND2X0 U6385 ( .IN1(g3201), .IN2(n4329), .QN(n3702) );
  NAND4X0 U6386 ( .IN1(g785), .IN2(g789), .IN3(n4047), .IN4(n4048), .QN(n3228)
         );
  NOR2X0 U6387 ( .IN1(n4391), .IN2(n4321), .QN(n4047) );
  NOR4X0 U6388 ( .IN1(n4289), .IN2(n4567), .IN3(n4559), .IN4(n4327), .QN(n4048) );
  NAND4X0 U6389 ( .IN1(g97), .IN2(g101), .IN3(n4052), .IN4(n4053), .QN(n3239)
         );
  NOR2X0 U6390 ( .IN1(n4392), .IN2(n4322), .QN(n4052) );
  NOR4X0 U6391 ( .IN1(n4290), .IN2(n4569), .IN3(n4561), .IN4(n4328), .QN(n4053) );
  AO222X1 U6392 ( .IN1(g2486), .IN2(n4608), .IN3(test_so80), .IN4(n4606), 
        .IN5(g2483), .IN6(n4610), .Q(n3192) );
  AO222X1 U6393 ( .IN1(g1792), .IN2(n4620), .IN3(g1795), .IN4(n4618), .IN5(
        g1789), .IN6(n4622), .Q(n3208) );
  AO222X1 U6394 ( .IN1(g411), .IN2(n4641), .IN3(g414), .IN4(n4640), .IN5(g408), 
        .IN6(n4643), .Q(n3233) );
  AO222X1 U6395 ( .IN1(g1095), .IN2(g5472), .IN3(g1101), .IN4(n4630), .IN5(
        g1098), .IN6(g6712), .Q(n3221) );
  NOR2X0 U6396 ( .IN1(n3706), .IN2(g3201), .QN(n3932) );
  NAND2X0 U6397 ( .IN1(n3945), .IN2(n3946), .QN(g25489) );
  NAND2X0 U6398 ( .IN1(n3947), .IN2(n4333), .QN(n3945) );
  NAND4X0 U6399 ( .IN1(g3142), .IN2(g3097), .IN3(g3151), .IN4(n3947), .QN(
        n3946) );
  AO221X1 U6400 ( .IN1(n3948), .IN2(n4424), .IN3(n3935), .IN4(n4301), .IN5(
        test_so10), .Q(n3947) );
  NOR2X0 U6401 ( .IN1(n4329), .IN2(g3188), .QN(n3933) );
  OA222X1 U6402 ( .IN1(n4524), .IN2(g2479), .IN3(n4509), .IN4(test_so82), 
        .IN5(n4516), .IN6(g2478), .Q(n2967) );
  OA222X1 U6403 ( .IN1(n4525), .IN2(g1785), .IN3(n4511), .IN4(g1783), .IN5(
        n4518), .IN6(test_so60), .Q(n2971) );
  OA222X1 U6404 ( .IN1(n4673), .IN2(g1090), .IN3(n4669), .IN4(g1089), .IN5(
        n4671), .IN6(g1091), .Q(n2975) );
  OA222X1 U6405 ( .IN1(n4676), .IN2(g404), .IN3(n4506), .IN4(g402), .IN5(n4520), .IN6(g403), .Q(n2978) );
  NAND2X0 U6406 ( .IN1(g3204), .IN2(n3938), .QN(n3706) );
  NAND2X0 U6407 ( .IN1(n3199), .IN2(g2257), .QN(n2791) );
  NAND2X0 U6408 ( .IN1(n3215), .IN2(g1563), .QN(n2610) );
  NAND2X0 U6409 ( .IN1(n3229), .IN2(g869), .QN(n2631) );
  NAND2X0 U6410 ( .IN1(n3240), .IN2(g181), .QN(n2651) );
  NAND2X0 U6411 ( .IN1(g2703), .IN2(n4426), .QN(n4186) );
  NAND2X0 U6412 ( .IN1(g2009), .IN2(n4427), .QN(n4189) );
  NAND2X0 U6413 ( .IN1(g1315), .IN2(n4428), .QN(n4192) );
  NAND2X0 U6414 ( .IN1(g629), .IN2(n4429), .QN(n4135) );
  NAND2X0 U6415 ( .IN1(DFF_16_n1), .IN2(DFF_15_n1), .QN(n3935) );
  NAND2X0 U6416 ( .IN1(g2707), .IN2(n4185), .QN(n4106) );
  NAND2X0 U6417 ( .IN1(g2013), .IN2(n4188), .QN(n4109) );
  NAND2X0 U6418 ( .IN1(g1319), .IN2(n4191), .QN(n4112) );
  NAND2X0 U6419 ( .IN1(g633), .IN2(n4134), .QN(n4115) );
  AO22X1 U6420 ( .IN1(n3447), .IN2(n4385), .IN3(n3449), .IN4(test_so79), .Q(
        n3710) );
  AO22X1 U6421 ( .IN1(n3459), .IN2(n4386), .IN3(n3461), .IN4(g1690), .Q(n3715)
         );
  AO22X1 U6422 ( .IN1(n3471), .IN2(n4387), .IN3(n3473), .IN4(g996), .Q(n3721)
         );
  AO22X1 U6423 ( .IN1(n3480), .IN2(n4388), .IN3(n3482), .IN4(g309), .Q(n3727)
         );
  AO222X1 U6424 ( .IN1(g617), .IN2(n4636), .IN3(test_so26), .IN4(n4633), .IN5(
        g614), .IN6(g6485), .Q(n2437) );
  AO222X1 U6425 ( .IN1(g608), .IN2(n4636), .IN3(g611), .IN4(n4634), .IN5(g605), 
        .IN6(n4638), .Q(n2432) );
  AO222X1 U6426 ( .IN1(g2691), .IN2(n4602), .IN3(g2694), .IN4(n4599), .IN5(
        g2688), .IN6(n4604), .Q(n2358) );
  AO222X1 U6427 ( .IN1(g1997), .IN2(n4614), .IN3(g2000), .IN4(n4611), .IN5(
        g1994), .IN6(n4616), .Q(n2286) );
  AO222X1 U6428 ( .IN1(g1303), .IN2(n4626), .IN3(g1306), .IN4(n4623), .IN5(
        g1300), .IN6(n4628), .Q(n2214) );
  AO222X1 U6429 ( .IN1(test_so90), .IN2(n4602), .IN3(g2685), .IN4(n4600), 
        .IN5(g2679), .IN6(g7302), .Q(n2353) );
  AO222X1 U6430 ( .IN1(g1988), .IN2(n4614), .IN3(g1991), .IN4(n4612), .IN5(
        g1985), .IN6(g7052), .Q(n2281) );
  AO222X1 U6431 ( .IN1(g1294), .IN2(n4626), .IN3(g1297), .IN4(n4624), .IN5(
        g1291), .IN6(g6750), .Q(n2209) );
  AND3X1 U6432 ( .IN1(n2397), .IN2(n3955), .IN3(n3956), .Q(n3949) );
  OR2X1 U6433 ( .IN1(n4306), .IN2(g2803), .Q(n3955) );
  OA222X1 U6434 ( .IN1(g2804), .IN2(n4356), .IN3(g2802), .IN4(n4292), .IN5(
        n3957), .IN6(n3958), .Q(n3956) );
  NAND4X0 U6435 ( .IN1(n3959), .IN2(n3960), .IN3(n3961), .IN4(n3962), .QN(
        n3958) );
  AND3X1 U6436 ( .IN1(n2325), .IN2(n3975), .IN3(n3976), .Q(n3952) );
  OR2X1 U6437 ( .IN1(n4307), .IN2(g2109), .Q(n3975) );
  OA222X1 U6438 ( .IN1(g2110), .IN2(n4357), .IN3(g2108), .IN4(n4293), .IN5(
        n3977), .IN6(n3978), .Q(n3976) );
  NAND4X0 U6439 ( .IN1(n3979), .IN2(n3980), .IN3(n3981), .IN4(n3982), .QN(
        n3978) );
  AND3X1 U6440 ( .IN1(n2253), .IN2(n3997), .IN3(n3998), .Q(n3972) );
  OR2X1 U6441 ( .IN1(n4308), .IN2(g1415), .Q(n3997) );
  OA222X1 U6442 ( .IN1(g1416), .IN2(n4358), .IN3(test_so51), .IN4(n4294), 
        .IN5(n3999), .IN6(n4000), .Q(n3998) );
  NAND4X0 U6443 ( .IN1(n4001), .IN2(n4002), .IN3(n4003), .IN4(n4004), .QN(
        n4000) );
  AND3X1 U6444 ( .IN1(n2475), .IN2(n4015), .IN3(n4016), .Q(n3992) );
  OR2X1 U6445 ( .IN1(n4309), .IN2(g729), .Q(n4015) );
  OA222X1 U6446 ( .IN1(g730), .IN2(n4359), .IN3(g728), .IN4(n4295), .IN5(n4017), .IN6(n4018), .Q(n4016) );
  NAND4X0 U6447 ( .IN1(n4019), .IN2(n4020), .IN3(n4021), .IN4(n4022), .QN(
        n4018) );
  OA222X1 U6448 ( .IN1(n3902), .IN2(n4343), .IN3(n3708), .IN4(n3695), .IN5(
        n3903), .IN6(n4447), .Q(n3923) );
  OA222X1 U6449 ( .IN1(n3902), .IN2(n4344), .IN3(n1626), .IN4(n3695), .IN5(
        n3903), .IN6(n4448), .Q(n3931) );
  OA221X1 U6450 ( .IN1(n3912), .IN2(n4445), .IN3(n3913), .IN4(n4340), .IN5(
        n3941), .Q(n3928) );
  OA222X1 U6451 ( .IN1(n3699), .IN2(n4332), .IN3(n3915), .IN4(n4446), .IN5(
        n3703), .IN6(n4301), .Q(n3941) );
  NAND2X0 U6452 ( .IN1(g2746), .IN2(n3746), .QN(n3681) );
  NAND2X0 U6453 ( .IN1(g2720), .IN2(n4105), .QN(n3747) );
  NAND2X0 U6454 ( .IN1(g2052), .IN2(n3754), .QN(n3489) );
  NAND2X0 U6455 ( .IN1(g2026), .IN2(n4108), .QN(n3755) );
  NAND2X0 U6456 ( .IN1(g1358), .IN2(n3784), .QN(n3493) );
  NAND2X0 U6457 ( .IN1(g1332), .IN2(n4111), .QN(n3785) );
  NAND2X0 U6458 ( .IN1(g672), .IN2(n3814), .QN(n3497) );
  NAND2X0 U6459 ( .IN1(g646), .IN2(n4114), .QN(n3815) );
  ISOLANDX1 U6460 ( .D(g3233), .ISO(g3230), .Q(n3700) );
  NOR2X0 U6461 ( .IN1(n4573), .IN2(n3198), .QN(n3449) );
  OA222X1 U6462 ( .IN1(n4324), .IN2(g2254), .IN3(n4682), .IN4(g2255), .IN5(
        n4367), .IN6(g2253), .Q(n4573) );
  NOR2X0 U6463 ( .IN1(n4574), .IN2(n3214), .QN(n3461) );
  OA222X1 U6464 ( .IN1(n4688), .IN2(g1560), .IN3(n4686), .IN4(g1561), .IN5(
        n4368), .IN6(g1559), .Q(n4574) );
  NOR2X0 U6465 ( .IN1(n4575), .IN2(n3228), .QN(n3473) );
  OA222X1 U6466 ( .IN1(n4323), .IN2(g866), .IN3(n4312), .IN4(g867), .IN5(n4691), .IN6(g865), .Q(n4575) );
  NOR2X0 U6467 ( .IN1(n4576), .IN2(n3239), .QN(n3482) );
  OA222X1 U6468 ( .IN1(n4698), .IN2(g178), .IN3(n4696), .IN4(g179), .IN5(n4369), .IN6(g177), .Q(n4576) );
  NAND4X0 U6469 ( .IN1(n4649), .IN2(g2908), .IN3(n4182), .IN4(n4183), .QN(
        n2483) );
  ISOLANDX1 U6470 ( .D(g2892), .ISO(n4305), .Q(n4182) );
  AND4X1 U6471 ( .IN1(n4291), .IN2(n4431), .IN3(n4330), .IN4(g2888), .Q(n4183)
         );
  NOR3X0 U6472 ( .IN1(g3201), .IN2(g3207), .IN3(g3188), .QN(n3934) );
  AND3X1 U6473 ( .IN1(DFF_132_n1), .IN2(DFF_134_n1), .IN3(DFF_131_n1), .Q(
        n3944) );
  NAND2X0 U6474 ( .IN1(g2753), .IN2(n3680), .QN(n3415) );
  NAND2X0 U6475 ( .IN1(g2059), .IN2(n3488), .QN(n3418) );
  NAND2X0 U6476 ( .IN1(g1365), .IN2(n3492), .QN(n3421) );
  NAND2X0 U6477 ( .IN1(g679), .IN2(n3496), .QN(n3243) );
  AND2X1 U6478 ( .IN1(n4073), .IN2(g3204), .Q(n3942) );
  NOR2X0 U6479 ( .IN1(g3036), .IN2(g3032), .QN(n4207) );
  INVX0 U6480 ( .IN(n4730), .QN(n4726) );
  INVX0 U6481 ( .IN(g2879), .QN(n4730) );
  NAND4X0 U6482 ( .IN1(n3694), .IN2(n3695), .IN3(n3696), .IN4(n3697), .QN(
        g27380) );
  NAND3X0 U6483 ( .IN1(n1748), .IN2(n1747), .IN3(n3707), .QN(n3694) );
  OA22X1_S38584 U6484 ( .IN1(n3701), .IN2(n3702), .IN3(n3703), .IN4(n4424), .Q(n3696)
         );
  OA221X1 U6485 ( .IN1(g3133), .IN2(n3698), .IN3(n3699), .IN4(n4425), .IN5(
        n3700), .Q(n3697) );
  INVX0 U6486 ( .IN(g3229), .QN(n4776) );
  OA221X1 U6487 ( .IN1(n3907), .IN2(n4442), .IN3(n3908), .IN4(n4341), .IN5(
        n3909), .Q(n3900) );
  OA22X1_S38584 U6488 ( .IN1(n3910), .IN2(n4345), .IN3(n3911), .IN4(n4450), .Q(n3909)
         );
  AO22X1 U6489 ( .IN1(DFF_328_n1), .IN2(n4430), .IN3(n4210), .IN4(g305), .Q(
        g21346) );
  NOR2X0 U6490 ( .IN1(n4641), .IN2(n4430), .QN(n4210) );
  OA221X1 U6491 ( .IN1(n3912), .IN2(n4443), .IN3(n3913), .IN4(n4342), .IN5(
        n3925), .Q(n3920) );
  OA222X1 U6492 ( .IN1(n3699), .IN2(DFF_155_n1), .IN3(n3915), .IN4(n4433), 
        .IN5(n3703), .IN6(n4333), .Q(n3925) );
  AND3X1 U6493 ( .IN1(n3160), .IN2(n3157), .IN3(n3423), .Q(g28148) );
  AND3X1 U6494 ( .IN1(n4522), .IN2(n3157), .IN3(n3682), .Q(g27131) );
  AND3X1 U6495 ( .IN1(n4526), .IN2(n3157), .IN3(n3886), .Q(g25940) );
  AND3X1 U6496 ( .IN1(n3164), .IN2(n3161), .IN3(n3426), .Q(g28147) );
  AND3X1 U6497 ( .IN1(n4523), .IN2(n3161), .IN3(n3685), .Q(g27129) );
  AND3X1 U6498 ( .IN1(n4527), .IN2(n3161), .IN3(n3889), .Q(g25938) );
  AND3X1 U6499 ( .IN1(n3168), .IN2(n3165), .IN3(n3429), .Q(g28146) );
  AND3X1 U6500 ( .IN1(n3431), .IN2(n3165), .IN3(n3688), .Q(g27123) );
  AND3X1 U6501 ( .IN1(n3690), .IN2(n3165), .IN3(n3892), .Q(g25935) );
  AND3X1 U6502 ( .IN1(n3172), .IN2(n3169), .IN3(n3432), .Q(g28145) );
  AND3X1 U6503 ( .IN1(n4521), .IN2(n3169), .IN3(n3691), .Q(g27120) );
  AND3X1 U6504 ( .IN1(n4528), .IN2(n3169), .IN3(n3895), .Q(g25932) );
  AND3X1 U6505 ( .IN1(n3681), .IN2(n3678), .IN3(n3745), .Q(g26677) );
  OR2X1 U6506 ( .IN1(n3746), .IN2(g2746), .Q(n3745) );
  AND3X1 U6507 ( .IN1(n3489), .IN2(n3486), .IN3(n3753), .Q(g26671) );
  OR2X1 U6508 ( .IN1(n3754), .IN2(g2052), .Q(n3753) );
  AND3X1 U6509 ( .IN1(n3493), .IN2(n3490), .IN3(n3783), .Q(g26666) );
  OR2X1 U6510 ( .IN1(n3784), .IN2(g1358), .Q(n3783) );
  AND3X1 U6511 ( .IN1(n3497), .IN2(n3494), .IN3(n3813), .Q(g26660) );
  OR2X1 U6512 ( .IN1(n3814), .IN2(g672), .Q(n3813) );
  AND3X1 U6513 ( .IN1(n3415), .IN2(n3678), .IN3(n3679), .Q(g27243) );
  OR2X1 U6514 ( .IN1(n3680), .IN2(g2753), .Q(n3679) );
  AND3X1 U6515 ( .IN1(n3418), .IN2(n3486), .IN3(n3487), .Q(g27682) );
  OR2X1 U6516 ( .IN1(n3488), .IN2(g2059), .Q(n3487) );
  AND3X1 U6517 ( .IN1(n3421), .IN2(n3490), .IN3(n3491), .Q(g27678) );
  OR2X1 U6518 ( .IN1(n3492), .IN2(g1365), .Q(n3491) );
  AND3X1 U6519 ( .IN1(n3243), .IN2(n3494), .IN3(n3495), .Q(g27672) );
  OR2X1 U6520 ( .IN1(n3496), .IN2(g679), .Q(n3495) );
  AO22X1 U6521 ( .IN1(g2543), .IN2(n4455), .IN3(g8167), .IN4(n2097), .Q(g24237) );
  AO22X1 U6522 ( .IN1(g2540), .IN2(n4456), .IN3(g8087), .IN4(n2097), .Q(g24225) );
  AO22X1 U6523 ( .IN1(g2559), .IN2(n4455), .IN3(g8167), .IN4(n2109), .Q(g23047) );
  AO22X1 U6524 ( .IN1(g2555), .IN2(n4456), .IN3(g8087), .IN4(n2109), .Q(g23132) );
  AO22X1 U6525 ( .IN1(g2553), .IN2(n4455), .IN3(g8167), .IN4(n2096), .Q(g24226) );
  AO22X1 U6526 ( .IN1(g2552), .IN2(n4456), .IN3(g8087), .IN4(n2096), .Q(g24214) );
  AO22X1 U6527 ( .IN1(g2562), .IN2(n4455), .IN3(g8167), .IN4(n3448), .Q(g23133) );
  AO22X1 U6528 ( .IN1(g2561), .IN2(n4456), .IN3(g8087), .IN4(n3448), .Q(g23114) );
  AO22X1 U6529 ( .IN1(g1849), .IN2(n4457), .IN3(g8082), .IN4(n1995), .Q(g24230) );
  AO22X1 U6530 ( .IN1(g1846), .IN2(n4458), .IN3(g8012), .IN4(n1995), .Q(g24218) );
  AO22X1 U6531 ( .IN1(g1865), .IN2(n4457), .IN3(g8082), .IN4(n2008), .Q(g23030) );
  AO22X1 U6532 ( .IN1(g1861), .IN2(n4458), .IN3(g8012), .IN4(n2008), .Q(g23123) );
  AO22X1 U6533 ( .IN1(g1859), .IN2(n4457), .IN3(g8082), .IN4(n1994), .Q(g24219) );
  AO22X1 U6534 ( .IN1(g1858), .IN2(n4458), .IN3(g8012), .IN4(n1994), .Q(g24208) );
  AO22X1 U6535 ( .IN1(g1868), .IN2(n4457), .IN3(g8082), .IN4(n3460), .Q(g23124) );
  AO22X1 U6536 ( .IN1(g1867), .IN2(n4458), .IN3(g8012), .IN4(n3460), .Q(g23097) );
  AO22X1 U6537 ( .IN1(g1155), .IN2(n4459), .IN3(g8007), .IN4(n1893), .Q(g24222) );
  AO22X1 U6538 ( .IN1(g1152), .IN2(n4460), .IN3(g7961), .IN4(n1893), .Q(g24212) );
  AO22X1 U6539 ( .IN1(g1171), .IN2(n4459), .IN3(g8007), .IN4(n1906), .Q(g23014) );
  AO22X1 U6540 ( .IN1(g1167), .IN2(n4460), .IN3(g7961), .IN4(n1906), .Q(g23110) );
  AO22X1 U6541 ( .IN1(g1165), .IN2(n4459), .IN3(g8007), .IN4(n1892), .Q(g24213) );
  AO22X1 U6542 ( .IN1(g1164), .IN2(n4460), .IN3(g7961), .IN4(n1892), .Q(g24181) );
  AO22X1 U6543 ( .IN1(test_so44), .IN2(n4459), .IN3(g8007), .IN4(n3472), .Q(
        g23111) );
  AO22X1 U6544 ( .IN1(g1173), .IN2(n4460), .IN3(g7961), .IN4(n3472), .Q(g23081) );
  AO22X1 U6545 ( .IN1(test_so24), .IN2(n4461), .IN3(g7956), .IN4(n1789), .Q(
        g24215) );
  AO22X1 U6546 ( .IN1(g465), .IN2(n4462), .IN3(g7909), .IN4(n1789), .Q(g24206)
         );
  AO22X1 U6547 ( .IN1(g484), .IN2(n4461), .IN3(g7956), .IN4(n1802), .Q(g23000)
         );
  AO22X1 U6548 ( .IN1(g480), .IN2(n4462), .IN3(g7909), .IN4(n1802), .Q(g23092)
         );
  AO22X1 U6549 ( .IN1(g478), .IN2(n4461), .IN3(g7956), .IN4(n1788), .Q(g24207)
         );
  AO22X1 U6550 ( .IN1(g477), .IN2(n4462), .IN3(g7909), .IN4(n1788), .Q(g24178)
         );
  AO22X1 U6551 ( .IN1(g487), .IN2(n4461), .IN3(g7956), .IN4(n3481), .Q(g23093)
         );
  AO22X1 U6552 ( .IN1(g486), .IN2(n4462), .IN3(g7909), .IN4(n3481), .Q(g23067)
         );
  NAND2X0 U6553 ( .IN1(g2917), .IN2(n2484), .QN(n4099) );
  AO22X1 U6554 ( .IN1(g2533), .IN2(n4455), .IN3(n2092), .IN4(g8167), .Q(g23418) );
  AO22X1 U6555 ( .IN1(g2530), .IN2(n4456), .IN3(n2092), .IN4(g8087), .Q(g23407) );
  AO22X1 U6556 ( .IN1(test_so65), .IN2(n4457), .IN3(n1990), .IN4(g8082), .Q(
        g23413) );
  AO22X1 U6557 ( .IN1(g1836), .IN2(n4458), .IN3(n1990), .IN4(g8012), .Q(g23400) );
  AO22X1 U6558 ( .IN1(g1145), .IN2(n4459), .IN3(n1888), .IN4(g8007), .Q(g23406) );
  AO22X1 U6559 ( .IN1(g1142), .IN2(n4460), .IN3(n1888), .IN4(g7961), .Q(g23392) );
  AO22X1 U6560 ( .IN1(g458), .IN2(n4461), .IN3(n1784), .IN4(g7956), .Q(g23399)
         );
  AO22X1 U6561 ( .IN1(g455), .IN2(n4462), .IN3(n1784), .IN4(g7909), .Q(g23385)
         );
  ISOLANDX1 U6562 ( .D(n3938), .ISO(g3204), .Q(n3939) );
  ISOLANDX1 U6563 ( .D(n4073), .ISO(g3204), .Q(n3705) );
  NOR2X0 U6564 ( .IN1(n4577), .IN2(n4578), .QN(n3708) );
  AO22X1 U6565 ( .IN1(g2546), .IN2(n4463), .IN3(g2560), .IN4(n2097), .Q(g24250) );
  AO22X1 U6566 ( .IN1(g1852), .IN2(n4464), .IN3(g1866), .IN4(n1995), .Q(g24243) );
  AO22X1 U6567 ( .IN1(g1158), .IN2(n4465), .IN3(g1172), .IN4(n1893), .Q(g24235) );
  AO22X1 U6568 ( .IN1(g471), .IN2(n4466), .IN3(g485), .IN4(n1789), .Q(g24228)
         );
  AO22X1 U6569 ( .IN1(g2536), .IN2(n4463), .IN3(n2092), .IN4(g2560), .Q(g24209) );
  AO22X1 U6570 ( .IN1(g1842), .IN2(n4464), .IN3(n1990), .IN4(g1866), .Q(g24182) );
  AO22X1 U6571 ( .IN1(g1148), .IN2(n4465), .IN3(n1888), .IN4(g1172), .Q(g24179) );
  AO22X1 U6572 ( .IN1(g461), .IN2(n4466), .IN3(n1784), .IN4(g485), .Q(g24174)
         );
  AO22X1 U6573 ( .IN1(g3102), .IN2(n4494), .IN3(n4644), .IN4(n1817), .Q(g28425) );
  AO22X1 U6574 ( .IN1(test_so7), .IN2(n4383), .IN3(n4646), .IN4(n1817), .Q(
        g28421) );
  AO22X1 U6575 ( .IN1(g3100), .IN2(n4382), .IN3(n4648), .IN4(n1817), .Q(g28420) );
  AO22X1 U6576 ( .IN1(g2554), .IN2(n4463), .IN3(g2560), .IN4(n2096), .Q(g24238) );
  AO22X1 U6577 ( .IN1(g1860), .IN2(n4464), .IN3(g1866), .IN4(n1994), .Q(g24231) );
  AO22X1 U6578 ( .IN1(g1166), .IN2(n4465), .IN3(g1172), .IN4(n1892), .Q(g24223) );
  AO22X1 U6579 ( .IN1(g479), .IN2(n4466), .IN3(g485), .IN4(n1788), .Q(g24216)
         );
  AO22X1 U6580 ( .IN1(g3105), .IN2(n4494), .IN3(n4644), .IN4(n1818), .Q(g29941) );
  AO22X1 U6581 ( .IN1(g3104), .IN2(n4383), .IN3(n4646), .IN4(n1818), .Q(g29939) );
  AO22X1 U6582 ( .IN1(g3103), .IN2(n4382), .IN3(g8106), .IN4(n1818), .Q(g29936) );
  AO22X1 U6583 ( .IN1(g2539), .IN2(n4463), .IN3(g2560), .IN4(n2109), .Q(g23076) );
  AO22X1 U6584 ( .IN1(test_so87), .IN2(n4463), .IN3(g2560), .IN4(n3448), .Q(
        g21970) );
  AO22X1 U6585 ( .IN1(g1845), .IN2(n4464), .IN3(g1866), .IN4(n2008), .Q(g23058) );
  AO22X1 U6586 ( .IN1(g1869), .IN2(n4464), .IN3(g1866), .IN4(n3460), .Q(g23137) );
  AO22X1 U6587 ( .IN1(g1151), .IN2(n4465), .IN3(g1172), .IN4(n1906), .Q(g23039) );
  AO22X1 U6588 ( .IN1(g1175), .IN2(n4465), .IN3(g1172), .IN4(n3472), .Q(g23126) );
  AO22X1 U6589 ( .IN1(g464), .IN2(n4466), .IN3(g485), .IN4(n1802), .Q(g23022)
         );
  AO22X1 U6590 ( .IN1(g488), .IN2(n4466), .IN3(g485), .IN4(n3481), .Q(g23117)
         );
  AO22X1 U6591 ( .IN1(g2963), .IN2(n4707), .IN3(g2165), .IN4(n4732), .Q(g18957) );
  AO22X1 U6592 ( .IN1(test_so2), .IN2(n4703), .IN3(g2170), .IN4(n4733), .Q(
        g18836) );
  AO22X1 U6593 ( .IN1(g2969), .IN2(n4704), .IN3(g2175), .IN4(n4733), .Q(g18867) );
  AO22X1 U6594 ( .IN1(g2972), .IN2(n4706), .IN3(g2180), .IN4(n4732), .Q(g18906) );
  AO22X1 U6595 ( .IN1(g2975), .IN2(n4706), .IN3(g2185), .IN4(n4732), .Q(g18942) );
  AO22X1 U6596 ( .IN1(g2978), .IN2(n4707), .IN3(g2190), .IN4(n4732), .Q(g18968) );
  AO22X1 U6597 ( .IN1(g2981), .IN2(n4708), .IN3(g2195), .IN4(n4732), .Q(g18975) );
  AO22X1 U6598 ( .IN1(g2874), .IN2(n4705), .IN3(g2200), .IN4(n4732), .Q(g18885) );
  AO22X1 U6599 ( .IN1(g2935), .IN2(n4705), .IN3(g1471), .IN4(n4732), .Q(g18883) );
  AO22X1 U6600 ( .IN1(g2938), .IN2(n4704), .IN3(g1476), .IN4(n4733), .Q(g18866) );
  AO22X1 U6601 ( .IN1(g2941), .IN2(n4703), .IN3(g1481), .IN4(n4733), .Q(g18852) );
  AO22X1 U6602 ( .IN1(g2944), .IN2(n4702), .IN3(g1486), .IN4(n4733), .Q(g18835) );
  AO22X1 U6603 ( .IN1(g2947), .IN2(n4702), .IN3(g1491), .IN4(n4733), .Q(g18821) );
  AO22X1 U6604 ( .IN1(g2953), .IN2(n4701), .IN3(g1496), .IN4(n4733), .Q(g18803) );
  AO22X1 U6605 ( .IN1(g2956), .IN2(n4701), .IN3(g1501), .IN4(n4733), .Q(g18781) );
  AO22X1 U6606 ( .IN1(g2959), .IN2(n4700), .IN3(g1506), .IN4(n4733), .Q(g18754) );
  AO22X1 U6607 ( .IN1(g2380), .IN2(n4736), .IN3(n4757), .IN4(n4483), .Q(g24092) );
  AO22X1 U6608 ( .IN1(g1686), .IN2(n4736), .IN3(n4757), .IN4(n4484), .Q(g24083) );
  AO22X1 U6609 ( .IN1(g305), .IN2(n4736), .IN3(n4758), .IN4(n4485), .Q(g24059)
         );
  AO22X1 U6610 ( .IN1(g2516), .IN2(n4664), .IN3(n3709), .IN4(n4608), .Q(g26826) );
  AO22X1 U6611 ( .IN1(g2507), .IN2(n4664), .IN3(n4608), .IN4(n3710), .Q(g26822) );
  AO22X1 U6612 ( .IN1(g2495), .IN2(n4664), .IN3(n4608), .IN4(n2996), .Q(g29221) );
  AO22X1 U6613 ( .IN1(g2486), .IN2(n4664), .IN3(n4608), .IN4(n3180), .Q(g28773) );
  AO22X1 U6614 ( .IN1(g1822), .IN2(n4667), .IN3(n3711), .IN4(n4620), .Q(g26821) );
  AO22X1 U6615 ( .IN1(g1813), .IN2(n4667), .IN3(n4620), .IN4(n3715), .Q(g26815) );
  AO22X1 U6616 ( .IN1(g1801), .IN2(n4667), .IN3(n4620), .IN4(n2997), .Q(g29212) );
  AO22X1 U6617 ( .IN1(g1792), .IN2(n4667), .IN3(n4620), .IN4(n3188), .Q(g28760) );
  AO22X1 U6618 ( .IN1(g1128), .IN2(n4672), .IN3(n3716), .IN4(g6712), .Q(g26814) );
  AO22X1 U6619 ( .IN1(test_so38), .IN2(n4672), .IN3(g6712), .IN4(n3721), .Q(
        g26809) );
  AO22X1 U6620 ( .IN1(g1107), .IN2(n4672), .IN3(g6712), .IN4(n3005), .Q(g29204) );
  AO22X1 U6621 ( .IN1(g1098), .IN2(n4672), .IN3(g6712), .IN4(n3204), .Q(g28746) );
  AO22X1 U6622 ( .IN1(g2519), .IN2(n4663), .IN3(n3709), .IN4(n4606), .Q(g26827) );
  AO22X1 U6623 ( .IN1(g2513), .IN2(n4665), .IN3(n3709), .IN4(n4610), .Q(g26823) );
  AO22X1 U6624 ( .IN1(g2510), .IN2(n4663), .IN3(n4606), .IN4(n3710), .Q(g26825) );
  AO22X1 U6625 ( .IN1(g2504), .IN2(n4665), .IN3(n4610), .IN4(n3710), .Q(g26817) );
  AO22X1 U6626 ( .IN1(g2498), .IN2(n4663), .IN3(n4606), .IN4(n2996), .Q(g29226) );
  AO22X1 U6627 ( .IN1(g2492), .IN2(n4665), .IN3(n4610), .IN4(n2996), .Q(g29213) );
  AO22X1 U6628 ( .IN1(test_so80), .IN2(n4663), .IN3(n4606), .IN4(n3180), .Q(
        g28782) );
  AO22X1 U6629 ( .IN1(g2483), .IN2(n4665), .IN3(n4610), .IN4(n3180), .Q(g28763) );
  AO22X1 U6630 ( .IN1(test_so59), .IN2(n4666), .IN3(n3711), .IN4(n4618), .Q(
        g26824) );
  AO22X1 U6631 ( .IN1(g1819), .IN2(n4668), .IN3(n3711), .IN4(n4622), .Q(g26816) );
  AO22X1 U6632 ( .IN1(g1816), .IN2(n4666), .IN3(n4618), .IN4(n3715), .Q(g26820) );
  AO22X1 U6633 ( .IN1(g1810), .IN2(n4668), .IN3(n4622), .IN4(n3715), .Q(g26811) );
  AO22X1 U6634 ( .IN1(g1804), .IN2(n4666), .IN3(n4618), .IN4(n2997), .Q(g29218) );
  AO22X1 U6635 ( .IN1(g1798), .IN2(n4668), .IN3(n4622), .IN4(n2997), .Q(g29205) );
  AO22X1 U6636 ( .IN1(g1795), .IN2(n4666), .IN3(n4618), .IN4(n3188), .Q(g28771) );
  AO22X1 U6637 ( .IN1(g1789), .IN2(n4668), .IN3(n4622), .IN4(n3188), .Q(g28749) );
  AO22X1 U6638 ( .IN1(g1131), .IN2(n4670), .IN3(n3716), .IN4(n4630), .Q(g26818) );
  AO22X1 U6639 ( .IN1(g1125), .IN2(n4674), .IN3(n3716), .IN4(g5472), .Q(g26810) );
  AO22X1 U6640 ( .IN1(g1122), .IN2(n4670), .IN3(n4630), .IN4(n3721), .Q(g26813) );
  AO22X1 U6641 ( .IN1(g1116), .IN2(n4674), .IN3(g5472), .IN4(n3721), .Q(g26806) );
  AO22X1 U6642 ( .IN1(g1110), .IN2(n4670), .IN3(n4630), .IN4(n3005), .Q(g29209) );
  AO22X1 U6643 ( .IN1(g1104), .IN2(n4674), .IN3(g5472), .IN4(n3005), .Q(g29198) );
  AO22X1 U6644 ( .IN1(g1101), .IN2(n4670), .IN3(n4630), .IN4(n3204), .Q(g28758) );
  AO22X1 U6645 ( .IN1(g1095), .IN2(n4674), .IN3(g5472), .IN4(n3204), .Q(g28738) );
  AO22X1 U6646 ( .IN1(g444), .IN2(n4675), .IN3(n3722), .IN4(n4640), .Q(g26812)
         );
  AO22X1 U6647 ( .IN1(g441), .IN2(n4677), .IN3(n3722), .IN4(n4641), .Q(g26808)
         );
  AO22X1 U6648 ( .IN1(g438), .IN2(n4678), .IN3(n3722), .IN4(n4643), .Q(g26805)
         );
  AO22X1 U6649 ( .IN1(g435), .IN2(n4675), .IN3(n4640), .IN4(n3727), .Q(g26807)
         );
  AO22X1 U6650 ( .IN1(g432), .IN2(n4677), .IN3(n4641), .IN4(n3727), .Q(g26804)
         );
  AO22X1 U6651 ( .IN1(g429), .IN2(n4678), .IN3(n4643), .IN4(n3727), .Q(g26803)
         );
  AO22X1 U6652 ( .IN1(g423), .IN2(n4675), .IN3(n4640), .IN4(n3013), .Q(g29201)
         );
  AO22X1 U6653 ( .IN1(g420), .IN2(n4677), .IN3(n4641), .IN4(n3013), .Q(g29197)
         );
  AO22X1 U6654 ( .IN1(g417), .IN2(n4678), .IN3(n4643), .IN4(n3013), .Q(g29194)
         );
  AO22X1 U6655 ( .IN1(g414), .IN2(n4675), .IN3(n4640), .IN4(n3220), .Q(g28744)
         );
  AO22X1 U6656 ( .IN1(g411), .IN2(n4677), .IN3(n4641), .IN4(n3220), .Q(g28735)
         );
  AO22X1 U6657 ( .IN1(g408), .IN2(n4678), .IN3(n4643), .IN4(n3220), .Q(g28732)
         );
  AO22X1 U6658 ( .IN1(g2935), .IN2(n4731), .IN3(g4450), .IN4(n4713), .Q(g19178) );
  AO22X1 U6659 ( .IN1(g2938), .IN2(n4731), .IN3(g4200), .IN4(n4712), .Q(g19167) );
  AO22X1 U6660 ( .IN1(g2941), .IN2(n4732), .IN3(g3993), .IN4(n4710), .Q(g19157) );
  AO22X1 U6661 ( .IN1(g2944), .IN2(n4732), .IN3(g8175), .IN4(n4709), .Q(g19149) );
  AO22X1 U6662 ( .IN1(g2947), .IN2(n4732), .IN3(g8023), .IN4(n4708), .Q(g19144) );
  AO22X1 U6663 ( .IN1(g2953), .IN2(n4731), .IN3(g4321), .IN4(n4712), .Q(g19172) );
  AO22X1 U6664 ( .IN1(g2956), .IN2(n4732), .IN3(g4088), .IN4(n4711), .Q(g19162) );
  AO22X1 U6665 ( .IN1(g2959), .IN2(n4732), .IN3(g8249), .IN4(n4709), .Q(g19153) );
  AO22X1 U6666 ( .IN1(g2963), .IN2(n4731), .IN3(g7334), .IN4(n4716), .Q(g20417) );
  AO22X1 U6667 ( .IN1(test_so2), .IN2(n4731), .IN3(g6895), .IN4(n4715), .Q(
        g20376) );
  AO22X1 U6668 ( .IN1(g2969), .IN2(n4731), .IN3(g6442), .IN4(n4715), .Q(g20343) );
  AO22X1 U6669 ( .IN1(g2972), .IN2(n4731), .IN3(g6225), .IN4(n4714), .Q(g20310) );
  AO22X1 U6670 ( .IN1(g2975), .IN2(n4731), .IN3(g4590), .IN4(n4714), .Q(g19184) );
  AO22X1 U6671 ( .IN1(g2978), .IN2(n4731), .IN3(g4323), .IN4(n4713), .Q(g19173) );
  AO22X1 U6672 ( .IN1(g2981), .IN2(n4732), .IN3(g4090), .IN4(n4711), .Q(g19163) );
  AO22X1 U6673 ( .IN1(g2874), .IN2(n4732), .IN3(g8251), .IN4(n4710), .Q(g19154) );
  AO22X1 U6674 ( .IN1(g2565), .IN2(n4314), .IN3(n3841), .IN4(n4604), .Q(g26575) );
  AO22X1 U6675 ( .IN1(test_so68), .IN2(n4296), .IN3(n3842), .IN4(n4616), .Q(
        g26559) );
  AO22X1 U6676 ( .IN1(test_so47), .IN2(n4371), .IN3(n3844), .IN4(n4628), .Q(
        g26547) );
  AO22X1 U6677 ( .IN1(g490), .IN2(n4298), .IN3(n3846), .IN4(n4638), .Q(g26541)
         );
  AO22X1 U6678 ( .IN1(g2571), .IN2(n4299), .IN3(n3841), .IN4(n4600), .Q(g26616) );
  AO22X1 U6679 ( .IN1(g1877), .IN2(n4366), .IN3(n3842), .IN4(n4612), .Q(g26592) );
  AO22X1 U6680 ( .IN1(g1183), .IN2(n4300), .IN3(n3844), .IN4(n4624), .Q(g26569) );
  AO22X1 U6681 ( .IN1(g496), .IN2(n4313), .IN3(n3846), .IN4(n4634), .Q(g26553)
         );
  AO22X1 U6682 ( .IN1(n4754), .IN2(n4486), .IN3(g992), .IN4(n4736), .Q(g24072)
         );
  AO22X1 U6683 ( .IN1(g2568), .IN2(n4370), .IN3(n3841), .IN4(n4602), .Q(g26596) );
  AO22X1 U6684 ( .IN1(g1874), .IN2(n4315), .IN3(n3842), .IN4(n4614), .Q(g26573) );
  AO22X1 U6685 ( .IN1(g1180), .IN2(n4316), .IN3(n3844), .IN4(n4626), .Q(g26557) );
  AO22X1 U6686 ( .IN1(g493), .IN2(n4372), .IN3(n3846), .IN4(n4636), .Q(g26545)
         );
  AO22X1 U6687 ( .IN1(g3107), .IN2(n4383), .IN3(n4646), .IN4(g30072), .Q(
        g30798) );
  AO22X1 U6688 ( .IN1(g3106), .IN2(n4382), .IN3(n4648), .IN4(g30072), .Q(
        g30796) );
  AO22X1 U6689 ( .IN1(g3108), .IN2(n4494), .IN3(n4644), .IN4(g30072), .Q(
        g30801) );
  OA22X1_S38584 U6690 ( .IN1(n4735), .IN2(n4490), .IN3(n4746), .IN4(DFF_1503_n1), .Q(
        n2334) );
  OA22X1_S38584 U6691 ( .IN1(n4735), .IN2(n4491), .IN3(n4744), .IN4(DFF_1153_n1), .Q(
        n2262) );
  OA22X1_S38584 U6692 ( .IN1(n4489), .IN2(n4736), .IN3(n4745), .IN4(DFF_803_n1), .Q(
        n2190) );
  OA22X1_S38584 U6693 ( .IN1(n4742), .IN2(DFF_453_n1), .IN3(n4736), .IN4(n4492), .Q(
        n2406) );
  AOI21X1 U6694 ( .IN1(n4579), .IN2(g2580), .IN3(n4580), .QN(g30061) );
  AOI221X1 U6695 ( .IN1(g28990), .IN2(n4602), .IN3(g16437), .IN4(n4370), .IN5(
        g2580), .QN(n4580) );
  NAND2X0 U6696 ( .IN1(n3708), .IN2(g3142), .QN(n3948) );
  XOR2X1 U6697 ( .IN1(n3712), .IN2(n2110), .Q(n3709) );
  NAND3X0 U6698 ( .IN1(n3443), .IN2(n2101), .IN3(test_so79), .QN(n3712) );
  INVX0 U6699 ( .IN(n3444), .QN(n2101) );
  XOR2X1 U6700 ( .IN1(n3718), .IN2(n2007), .Q(n3711) );
  NAND3X0 U6701 ( .IN1(n3455), .IN2(n1999), .IN3(g1690), .QN(n3718) );
  INVX0 U6702 ( .IN(n3456), .QN(n1999) );
  XOR2X1 U6703 ( .IN1(n3724), .IN2(n1905), .Q(n3716) );
  NAND3X0 U6704 ( .IN1(n3467), .IN2(n1897), .IN3(g996), .QN(n3724) );
  INVX0 U6705 ( .IN(n3468), .QN(n1897) );
  XOR2X1 U6706 ( .IN1(n3729), .IN2(n1801), .Q(n3722) );
  NAND3X0 U6707 ( .IN1(n3476), .IN2(n1793), .IN3(g309), .QN(n3729) );
  INVX0 U6708 ( .IN(n3477), .QN(n1793) );
  XNOR2X1 U6709 ( .IN1(n4228), .IN2(n4229), .Q(n2420) );
  XOR3X1 U6710 ( .IN1(n4231), .IN2(g8263), .IN3(DFF_1628_n1), .Q(n4228) );
  XOR3X1 U6711 ( .IN1(DFF_1625_n1), .IN2(n4230), .IN3(DFF_1626_n1), .Q(n4229)
         );
  XOR2X1 U6712 ( .IN1(g8259), .IN2(g8264), .Q(n4231) );
  XNOR2X1 U6713 ( .IN1(n4224), .IN2(n4225), .Q(n2421) );
  XOR3X1 U6714 ( .IN1(n4227), .IN2(g8269), .IN3(DFF_1618_n1), .Q(n4224) );
  XOR3X1 U6715 ( .IN1(DFF_1616_n1), .IN2(n4226), .IN3(DFF_1617_n1), .Q(n4225)
         );
  XOR2X1 U6716 ( .IN1(g8271), .IN2(g8270), .Q(n4227) );
  AND2X1 U6717 ( .IN1(n3944), .IN2(g3197), .Q(n3938) );
  ISOLANDX1 U6718 ( .D(n3944), .ISO(g3197), .Q(n4073) );
  NAND3X0 U6719 ( .IN1(g3207), .IN2(g3201), .IN3(n3936), .QN(n3908) );
  NAND3X0 U6720 ( .IN1(g3207), .IN2(n4406), .IN3(n3936), .QN(n3913) );
  AO21X1 U6721 ( .IN1(g8021), .IN2(DFF_18_n1), .IN3(n4733), .Q(n4279) );
  NAND3X0 U6722 ( .IN1(g3188), .IN2(n4329), .IN3(n3932), .QN(n3902) );
  NAND3X0 U6723 ( .IN1(g3207), .IN2(g3188), .IN3(n3932), .QN(n3911) );
  NAND3X0 U6724 ( .IN1(test_so79), .IN2(n1687), .IN3(n2967), .QN(n3749) );
  NAND3X0 U6725 ( .IN1(test_so79), .IN2(n3443), .IN3(n3444), .QN(n3436) );
  NAND3X0 U6726 ( .IN1(g1690), .IN2(n1630), .IN3(n2971), .QN(n3751) );
  NAND3X0 U6727 ( .IN1(g1690), .IN2(n3455), .IN3(n3456), .QN(n3440) );
  NAND3X0 U6728 ( .IN1(g996), .IN2(n1649), .IN3(n2975), .QN(n3758) );
  NAND3X0 U6729 ( .IN1(g996), .IN2(n3467), .IN3(n3468), .QN(n3452) );
  NAND3X0 U6730 ( .IN1(g309), .IN2(n1668), .IN3(n2978), .QN(n3788) );
  NAND3X0 U6731 ( .IN1(g309), .IN2(n3476), .IN3(n3477), .QN(n3464) );
  OA22X1_S38584 U6732 ( .IN1(g2810), .IN2(n2146), .IN3(n3949), .IN4(n3951), .Q(g25280) );
  OA22X1_S38584 U6733 ( .IN1(g2809), .IN2(n2145), .IN3(n3949), .IN4(n3954), .Q(g25272) );
  OA22X1_S38584 U6734 ( .IN1(g2116), .IN2(n2044), .IN3(n3952), .IN4(n3971), .Q(g25271) );
  OA22X1_S38584 U6735 ( .IN1(g2115), .IN2(n2043), .IN3(n3952), .IN4(n3974), .Q(g25268) );
  OA22X1_S38584 U6736 ( .IN1(g1422), .IN2(n1942), .IN3(n3972), .IN4(n3991), .Q(g25267) );
  OA22X1_S38584 U6737 ( .IN1(g1421), .IN2(n1941), .IN3(n3972), .IN4(n3996), .Q(g25263) );
  OA22X1_S38584 U6738 ( .IN1(g736), .IN2(n1841), .IN3(n3992), .IN4(n4013), .Q(g25262)
         );
  OA22X1_S38584 U6739 ( .IN1(g735), .IN2(n1840), .IN3(n3992), .IN4(n4014), .Q(g25260)
         );
  AOI222X1 U6740 ( .IN1(g567), .IN2(n4636), .IN3(g489), .IN4(n4634), .IN5(g565), .IN6(n4638), .QN(g12457) );
  AOI222X1 U6741 ( .IN1(g571), .IN2(n4636), .IN3(g573), .IN4(n4634), .IN5(g569), .IN6(g6485), .QN(g12487) );
  AOI222X1 U6742 ( .IN1(g2641), .IN2(n4602), .IN3(g2564), .IN4(n4600), .IN5(
        g2639), .IN6(n4604), .QN(g12499) );
  AOI222X1 U6743 ( .IN1(g2645), .IN2(n4602), .IN3(g2647), .IN4(n4600), .IN5(
        g2643), .IN6(g7302), .QN(g12539) );
  AOI222X1 U6744 ( .IN1(g1947), .IN2(n4614), .IN3(g1870), .IN4(n4612), .IN5(
        g1945), .IN6(n4616), .QN(g12482) );
  AOI222X1 U6745 ( .IN1(g1951), .IN2(n4614), .IN3(g1953), .IN4(n4612), .IN5(
        g1949), .IN6(g7052), .QN(g12524) );
  AOI222X1 U6746 ( .IN1(g1253), .IN2(n4626), .IN3(g1176), .IN4(n4624), .IN5(
        g1251), .IN6(g6750), .QN(g12467) );
  AOI222X1 U6747 ( .IN1(g1257), .IN2(n4626), .IN3(g1259), .IN4(n4624), .IN5(
        g1255), .IN6(n4628), .QN(g12507) );
  NBUFFX2 U6748 ( .IN(g551), .Q(n4636) );
  OA22X1_S38584 U6749 ( .IN1(g2808), .IN2(n2147), .IN3(n3949), .IN4(n3950), .Q(g25288) );
  OA22X1_S38584 U6750 ( .IN1(g2114), .IN2(n2045), .IN3(n3952), .IN4(n3953), .Q(g25279) );
  OA22X1_S38584 U6751 ( .IN1(g1420), .IN2(n1943), .IN3(n3972), .IN4(n3973), .Q(g25270) );
  OA22X1_S38584 U6752 ( .IN1(g734), .IN2(n1842), .IN3(n3992), .IN4(n3993), .Q(g25266)
         );
  OA22X1_S38584 U6753 ( .IN1(n1577), .IN2(n4211), .IN3(g8096), .IN4(n4733), .Q(g20874) );
  INVX0 U6754 ( .IN(n4197), .QN(n1577) );
  NAND2X0 U6755 ( .IN1(n4198), .IN2(n4731), .QN(n4211) );
  OA22X1_S38584 U6756 ( .IN1(n1578), .IN2(n4199), .IN3(g7519), .IN4(n4733), .Q(g21878) );
  INVX0 U6757 ( .IN(n4194), .QN(n1578) );
  NAND2X0 U6758 ( .IN1(n4195), .IN2(n4731), .QN(n4199) );
  NBUFFX2 U6759 ( .IN(g2625), .Q(n4602) );
  NBUFFX2 U6760 ( .IN(g1931), .Q(n4614) );
  NBUFFX2 U6761 ( .IN(g1237), .Q(n4626) );
  OA22X1_S38584 U6762 ( .IN1(g2235), .IN2(n2088), .IN3(n3062), .IN4(n4169), .Q(g22184) );
  OA22X1_S38584 U6763 ( .IN1(g2237), .IN2(n2086), .IN3(n3062), .IN4(n4170), .Q(g22172) );
  OA22X1_S38584 U6764 ( .IN1(g2236), .IN2(n2084), .IN3(n3062), .IN4(n4172), .Q(g22155) );
  OA22X1_S38584 U6765 ( .IN1(g1541), .IN2(n1986), .IN3(n3094), .IN4(n4171), .Q(g22168) );
  OA22X1_S38584 U6766 ( .IN1(g1543), .IN2(n1984), .IN3(n3094), .IN4(n4173), .Q(g22151) );
  OA22X1_S38584 U6767 ( .IN1(g1542), .IN2(n1982), .IN3(n3094), .IN4(n4175), .Q(g22132) );
  OA22X1_S38584 U6768 ( .IN1(g159), .IN2(n1780), .IN3(n3154), .IN4(n4177), .Q(g22124)
         );
  OA22X1_S38584 U6769 ( .IN1(g161), .IN2(n1778), .IN3(n3154), .IN4(n4179), .Q(g22102)
         );
  OA22X1_S38584 U6770 ( .IN1(g160), .IN2(n1776), .IN3(n3154), .IN4(n4180), .Q(g22081)
         );
  OA22X1_S38584 U6771 ( .IN1(g2238), .IN2(n2088), .IN3(n2666), .IN4(n4169), .Q(g22194) );
  OA22X1_S38584 U6772 ( .IN1(test_so75), .IN2(n2086), .IN3(n2666), .IN4(n4170), .Q(
        g22185) );
  OA22X1_S38584 U6773 ( .IN1(g2239), .IN2(n2084), .IN3(n2666), .IN4(n4172), .Q(g22173) );
  OA22X1_S38584 U6774 ( .IN1(g2232), .IN2(n2088), .IN3(n4287), .IN4(n4169), .Q(g22171) );
  OA22X1_S38584 U6775 ( .IN1(g2229), .IN2(n2088), .IN3(n4563), .IN4(n4169), .Q(g22153) );
  OA22X1_S38584 U6776 ( .IN1(g2226), .IN2(n2088), .IN3(n4555), .IN4(n4169), .Q(g22138) );
  OA22X1_S38584 U6777 ( .IN1(g2223), .IN2(n2088), .IN3(n4325), .IN4(n4169), .Q(g22115) );
  OA22X1_S38584 U6778 ( .IN1(g2220), .IN2(n2088), .IN3(n4389), .IN4(n4169), .Q(g22097) );
  OA22X1_S38584 U6779 ( .IN1(g2217), .IN2(n2088), .IN3(n4319), .IN4(n4169), .Q(g22076) );
  OA22X1_S38584 U6780 ( .IN1(g2208), .IN2(n2088), .IN3(n4373), .IN4(n4169), .Q(g22200) );
  OA22X1_S38584 U6781 ( .IN1(g2205), .IN2(n2088), .IN3(n4377), .IN4(n4169), .Q(g22192) );
  OA22X1_S38584 U6782 ( .IN1(g1544), .IN2(n1986), .IN3(n2681), .IN4(n4171), .Q(g22180) );
  OA22X1_S38584 U6783 ( .IN1(g1546), .IN2(n1984), .IN3(n2681), .IN4(n4173), .Q(g22169) );
  OA22X1_S38584 U6784 ( .IN1(g1545), .IN2(n1982), .IN3(n2681), .IN4(n4175), .Q(g22152) );
  OA22X1_S38584 U6785 ( .IN1(g1538), .IN2(n1986), .IN3(n4288), .IN4(n4171), .Q(g22150) );
  OA22X1_S38584 U6786 ( .IN1(g1535), .IN2(n1986), .IN3(n4565), .IN4(n4171), .Q(g22130) );
  OA22X1_S38584 U6787 ( .IN1(g1532), .IN2(n1986), .IN3(n4557), .IN4(n4171), .Q(g22112) );
  OA22X1_S38584 U6788 ( .IN1(g1529), .IN2(n1986), .IN3(n4326), .IN4(n4171), .Q(g22090) );
  OA22X1_S38584 U6789 ( .IN1(g1526), .IN2(n1986), .IN3(n4390), .IN4(n4171), .Q(g22073) );
  OA22X1_S38584 U6790 ( .IN1(g1523), .IN2(n1986), .IN3(n4320), .IN4(n4171), .Q(g22057) );
  OA22X1_S38584 U6791 ( .IN1(g1514), .IN2(n1986), .IN3(n4374), .IN4(n4171), .Q(g22191) );
  OA22X1_S38584 U6792 ( .IN1(g1511), .IN2(n1986), .IN3(n4378), .IN4(n4171), .Q(g22178) );
  OA22X1_S38584 U6793 ( .IN1(g850), .IN2(n1884), .IN3(n2696), .IN4(n4174), .Q(g22164)
         );
  OA22X1_S38584 U6794 ( .IN1(g852), .IN2(n1882), .IN3(n2696), .IN4(n4176), .Q(g22148)
         );
  OA22X1_S38584 U6795 ( .IN1(g851), .IN2(n1880), .IN3(n2696), .IN4(n4178), .Q(g22129)
         );
  OA22X1_S38584 U6796 ( .IN1(g847), .IN2(n1884), .IN3(n3227), .IN4(n4174), .Q(g22147)
         );
  OA22X1_S38584 U6797 ( .IN1(g849), .IN2(n1882), .IN3(n3227), .IN4(n4176), .Q(g22128)
         );
  OA22X1_S38584 U6798 ( .IN1(g848), .IN2(n1880), .IN3(n3227), .IN4(n4178), .Q(g22106)
         );
  OA22X1_S38584 U6799 ( .IN1(g844), .IN2(n1884), .IN3(n4289), .IN4(n4174), .Q(g22127)
         );
  OA22X1_S38584 U6800 ( .IN1(g841), .IN2(n1884), .IN3(n4567), .IN4(n4174), .Q(g22104)
         );
  OA22X1_S38584 U6801 ( .IN1(g838), .IN2(n1884), .IN3(n4559), .IN4(n4174), .Q(g22087)
         );
  OA22X1_S38584 U6802 ( .IN1(g835), .IN2(n1884), .IN3(n4327), .IN4(n4174), .Q(g22066)
         );
  OA22X1_S38584 U6803 ( .IN1(g832), .IN2(n1884), .IN3(n4391), .IN4(n4174), .Q(g22054)
         );
  OA22X1_S38584 U6804 ( .IN1(g829), .IN2(n1884), .IN3(n4321), .IN4(n4174), .Q(g22040)
         );
  OA22X1_S38584 U6805 ( .IN1(g820), .IN2(n1884), .IN3(n4375), .IN4(n4174), .Q(g22177)
         );
  OA22X1_S38584 U6806 ( .IN1(g817), .IN2(n1884), .IN3(n4379), .IN4(n4174), .Q(g22162)
         );
  OA22X1_S38584 U6807 ( .IN1(g162), .IN2(n1780), .IN3(n2714), .IN4(n4177), .Q(g22143)
         );
  OA22X1_S38584 U6808 ( .IN1(g164), .IN2(n1778), .IN3(n2714), .IN4(n4179), .Q(g22125)
         );
  OA22X1_S38584 U6809 ( .IN1(test_so12), .IN2(n1776), .IN3(n2714), .IN4(n4180), .Q(
        g22103) );
  OA22X1_S38584 U6810 ( .IN1(g156), .IN2(n1780), .IN3(n4290), .IN4(n4177), .Q(g22101)
         );
  OA22X1_S38584 U6811 ( .IN1(g153), .IN2(n1780), .IN3(n4569), .IN4(n4177), .Q(g22079)
         );
  OA22X1_S38584 U6812 ( .IN1(g150), .IN2(n1780), .IN3(n4561), .IN4(n4177), .Q(g22063)
         );
  OA22X1_S38584 U6813 ( .IN1(g147), .IN2(n1780), .IN3(n4328), .IN4(n4177), .Q(g22047)
         );
  OA22X1_S38584 U6814 ( .IN1(test_so11), .IN2(n1780), .IN3(n4392), .IN4(n4177), .Q(
        g22037) );
  OA22X1_S38584 U6815 ( .IN1(g141), .IN2(n1780), .IN3(n4322), .IN4(n4177), .Q(g22030)
         );
  OA22X1_S38584 U6816 ( .IN1(g132), .IN2(n1780), .IN3(n4376), .IN4(n4177), .Q(g22161)
         );
  OA22X1_S38584 U6817 ( .IN1(g129), .IN2(n1780), .IN3(n4380), .IN4(n4177), .Q(g22141)
         );
  OA22X1_S38584 U6818 ( .IN1(g2807), .IN2(n2164), .IN3(n2125), .IN4(n3678), .Q(g21047) );
  OA22X1_S38584 U6819 ( .IN1(g2804), .IN2(n2164), .IN3(n2126), .IN4(n3678), .Q(g21028) );
  OA22X1_S38584 U6820 ( .IN1(g2113), .IN2(n2062), .IN3(n2023), .IN4(n3486), .Q(g21023) );
  OA22X1_S38584 U6821 ( .IN1(g2110), .IN2(n2062), .IN3(n2024), .IN4(n3486), .Q(g21002) );
  OA22X1_S38584 U6822 ( .IN1(g1419), .IN2(n1960), .IN3(n1921), .IN4(n3490), .Q(g20997) );
  OA22X1_S38584 U6823 ( .IN1(g1416), .IN2(n1960), .IN3(n1922), .IN4(n3490), .Q(g20975) );
  OA22X1_S38584 U6824 ( .IN1(g733), .IN2(n1859), .IN3(n1819), .IN4(n3494), .Q(g20970)
         );
  OA22X1_S38584 U6825 ( .IN1(g730), .IN2(n1859), .IN3(n1820), .IN4(n3494), .Q(g20947)
         );
  OA22X1_S38584 U6826 ( .IN1(g2806), .IN2(n2162), .IN3(n2125), .IN4(n4153), .Q(g21029) );
  OA22X1_S38584 U6827 ( .IN1(g2803), .IN2(n2162), .IN3(n2126), .IN4(n4153), .Q(g21007) );
  OA22X1_S38584 U6828 ( .IN1(g2112), .IN2(n2060), .IN3(n2023), .IN4(n4159), .Q(g21003) );
  OA22X1_S38584 U6829 ( .IN1(g2109), .IN2(n2060), .IN3(n2024), .IN4(n4159), .Q(g20980) );
  OA22X1_S38584 U6830 ( .IN1(g1418), .IN2(n1958), .IN3(n1921), .IN4(n4165), .Q(g20976) );
  OA22X1_S38584 U6831 ( .IN1(g1415), .IN2(n1958), .IN3(n1922), .IN4(n4165), .Q(g20952) );
  OA22X1_S38584 U6832 ( .IN1(g732), .IN2(n1857), .IN3(n1819), .IN4(n4168), .Q(g20948)
         );
  OA22X1_S38584 U6833 ( .IN1(g729), .IN2(n1857), .IN3(n1820), .IN4(n4168), .Q(g20924)
         );
  NBUFFX2 U6834 ( .IN(g1092), .Q(g6712) );
  OA22X1_S38584 U6835 ( .IN1(n3915), .IN2(n4449), .IN3(n3699), .IN4(DFF_156_n1), .Q(
        n3914) );
  OA22X1_S38584 U6836 ( .IN1(n3910), .IN2(n4346), .IN3(n3911), .IN4(n4451), .Q(n3937)
         );
  OA22X1_S38584 U6837 ( .IN1(n3910), .IN2(n4347), .IN3(n3911), .IN4(n4452), .Q(n3924)
         );
  OA22X1_S38584 U6838 ( .IN1(n3905), .IN2(n4348), .IN3(n3906), .IN4(n4453), .Q(n3904)
         );
  OA22X1_S38584 U6839 ( .IN1(g2253), .IN2(n1590), .IN3(n3198), .IN4(n4031), .Q(g25259) );
  OA22X1_S38584 U6840 ( .IN1(g2255), .IN2(n1591), .IN3(n3198), .IN4(n4032), .Q(g25257) );
  OA22X1_S38584 U6841 ( .IN1(g2254), .IN2(n1593), .IN3(n3198), .IN4(n4034), .Q(g25253) );
  OA22X1_S38584 U6842 ( .IN1(g2250), .IN2(n1590), .IN3(n4377), .IN4(n4031), .Q(g25256) );
  OA22X1_S38584 U6843 ( .IN1(g2252), .IN2(n1591), .IN3(n4377), .IN4(n4032), .Q(g25252) );
  OA22X1_S38584 U6844 ( .IN1(g2251), .IN2(n1593), .IN3(n4377), .IN4(n4034), .Q(g25247) );
  OA22X1_S38584 U6845 ( .IN1(g2247), .IN2(n1590), .IN3(n4373), .IN4(n4031), .Q(g25251) );
  OA22X1_S38584 U6846 ( .IN1(g2249), .IN2(n1591), .IN3(n4373), .IN4(n4032), .Q(g25246) );
  OA22X1_S38584 U6847 ( .IN1(g2248), .IN2(n1593), .IN3(n4373), .IN4(n4034), .Q(g25237) );
  OA22X1_S38584 U6848 ( .IN1(g2244), .IN2(n1590), .IN3(n4039), .IN4(n4031), .Q(g25245) );
  OA22X1_S38584 U6849 ( .IN1(g2246), .IN2(n1591), .IN3(n4039), .IN4(n4032), .Q(g25236) );
  OA22X1_S38584 U6850 ( .IN1(g2245), .IN2(n1593), .IN3(n4039), .IN4(n4034), .Q(g25227) );
  OA22X1_S38584 U6851 ( .IN1(g1559), .IN2(n1592), .IN3(n3214), .IN4(n4033), .Q(g25255) );
  OA22X1_S38584 U6852 ( .IN1(g1561), .IN2(n1594), .IN3(n3214), .IN4(n4037), .Q(g25250) );
  OA22X1_S38584 U6853 ( .IN1(g1560), .IN2(n1596), .IN3(n3214), .IN4(n4040), .Q(g25244) );
  OA22X1_S38584 U6854 ( .IN1(g1556), .IN2(n1592), .IN3(n4378), .IN4(n4033), .Q(g25249) );
  OA22X1_S38584 U6855 ( .IN1(g1558), .IN2(n1594), .IN3(n4378), .IN4(n4037), .Q(g25243) );
  OA22X1_S38584 U6856 ( .IN1(g1557), .IN2(n1596), .IN3(n4378), .IN4(n4040), .Q(g25235) );
  OA22X1_S38584 U6857 ( .IN1(test_so54), .IN2(n1592), .IN3(n4374), .IN4(n4033), .Q(
        g25242) );
  OA22X1_S38584 U6858 ( .IN1(g1555), .IN2(n1594), .IN3(n4374), .IN4(n4037), .Q(g25234) );
  OA22X1_S38584 U6859 ( .IN1(g1554), .IN2(n1596), .IN3(n4374), .IN4(n4040), .Q(g25225) );
  OA22X1_S38584 U6860 ( .IN1(g1550), .IN2(n1592), .IN3(n4045), .IN4(n4033), .Q(g25233) );
  OA22X1_S38584 U6861 ( .IN1(g1552), .IN2(n1594), .IN3(n4045), .IN4(n4037), .Q(g25224) );
  OA22X1_S38584 U6862 ( .IN1(g1551), .IN2(n1596), .IN3(n4045), .IN4(n4040), .Q(g25217) );
  OA22X1_S38584 U6863 ( .IN1(g865), .IN2(n1595), .IN3(n3228), .IN4(n4038), .Q(g25248)
         );
  OA22X1_S38584 U6864 ( .IN1(g867), .IN2(n1597), .IN3(n3228), .IN4(n4043), .Q(g25241)
         );
  OA22X1_S38584 U6865 ( .IN1(g866), .IN2(n1599), .IN3(n3228), .IN4(n4046), .Q(g25232)
         );
  OA22X1_S38584 U6866 ( .IN1(g862), .IN2(n1595), .IN3(n4379), .IN4(n4038), .Q(g25240)
         );
  OA22X1_S38584 U6867 ( .IN1(g864), .IN2(n1597), .IN3(n4379), .IN4(n4043), .Q(g25231)
         );
  OA22X1_S38584 U6868 ( .IN1(g863), .IN2(n1599), .IN3(n4379), .IN4(n4046), .Q(g25223)
         );
  OA22X1_S38584 U6869 ( .IN1(g859), .IN2(n1595), .IN3(n4375), .IN4(n4038), .Q(g25230)
         );
  OA22X1_S38584 U6870 ( .IN1(g861), .IN2(n1597), .IN3(n4375), .IN4(n4043), .Q(g25222)
         );
  OA22X1_S38584 U6871 ( .IN1(g860), .IN2(n1599), .IN3(n4375), .IN4(n4046), .Q(g25215)
         );
  OA22X1_S38584 U6872 ( .IN1(g856), .IN2(n1595), .IN3(n4050), .IN4(n4038), .Q(g25221)
         );
  OA22X1_S38584 U6873 ( .IN1(test_so33), .IN2(n1597), .IN3(n4050), .IN4(n4043), .Q(
        g25214) );
  OA22X1_S38584 U6874 ( .IN1(g857), .IN2(n1599), .IN3(n4050), .IN4(n4046), .Q(g25209)
         );
  OA22X1_S38584 U6875 ( .IN1(g177), .IN2(n1598), .IN3(n3239), .IN4(n4044), .Q(g25239)
         );
  OA22X1_S38584 U6876 ( .IN1(g179), .IN2(n1600), .IN3(n3239), .IN4(n4049), .Q(g25229)
         );
  OA22X1_S38584 U6877 ( .IN1(g178), .IN2(n1601), .IN3(n3239), .IN4(n4051), .Q(g25220)
         );
  OA22X1_S38584 U6878 ( .IN1(g174), .IN2(n1598), .IN3(n4380), .IN4(n4044), .Q(g25228)
         );
  OA22X1_S38584 U6879 ( .IN1(g176), .IN2(n1600), .IN3(n4380), .IN4(n4049), .Q(g25219)
         );
  OA22X1_S38584 U6880 ( .IN1(g175), .IN2(n1601), .IN3(n4380), .IN4(n4051), .Q(g25213)
         );
  OA22X1_S38584 U6881 ( .IN1(g171), .IN2(n1598), .IN3(n4376), .IN4(n4044), .Q(g25218)
         );
  OA22X1_S38584 U6882 ( .IN1(g173), .IN2(n1600), .IN3(n4376), .IN4(n4049), .Q(g25212)
         );
  OA22X1_S38584 U6883 ( .IN1(g172), .IN2(n1601), .IN3(n4376), .IN4(n4051), .Q(g25207)
         );
  OA22X1_S38584 U6884 ( .IN1(g168), .IN2(n1598), .IN3(n4054), .IN4(n4044), .Q(g25211)
         );
  OA22X1_S38584 U6885 ( .IN1(g170), .IN2(n1600), .IN3(n4054), .IN4(n4049), .Q(g25206)
         );
  OA22X1_S38584 U6886 ( .IN1(g169), .IN2(n1601), .IN3(n4054), .IN4(n4051), .Q(g25204)
         );
  OA21X1 U6887 ( .IN1(n3698), .IN2(DFF_140_n1), .IN3(n3700), .Q(n3943) );
  OA21X1 U6888 ( .IN1(g3128), .IN2(n3698), .IN3(n3700), .Q(n3926) );
  OA21X1 U6889 ( .IN1(n3698), .IN2(DFF_142_n1), .IN3(n3700), .Q(n3918) );
  OA22X1_S38584 U6890 ( .IN1(g2805), .IN2(n2165), .IN3(n2125), .IN4(n4146), .Q(g21063) );
  OA22X1_S38584 U6891 ( .IN1(g2802), .IN2(n2165), .IN3(n2126), .IN4(n4146), .Q(g21046) );
  OA22X1_S38584 U6892 ( .IN1(g2111), .IN2(n2063), .IN3(n2023), .IN4(n4150), .Q(g21042) );
  OA22X1_S38584 U6893 ( .IN1(g2108), .IN2(n2063), .IN3(n2024), .IN4(n4150), .Q(g21022) );
  OA22X1_S38584 U6894 ( .IN1(g1417), .IN2(n1961), .IN3(n1921), .IN4(n4156), .Q(g21018) );
  OA22X1_S38584 U6895 ( .IN1(test_so51), .IN2(n1961), .IN3(n1922), .IN4(n4156), .Q(
        g20996) );
  OA22X1_S38584 U6896 ( .IN1(g731), .IN2(n1860), .IN3(n1819), .IN4(n4162), .Q(g20992)
         );
  OA22X1_S38584 U6897 ( .IN1(g728), .IN2(n1860), .IN3(n1820), .IN4(n4162), .Q(g20969)
         );
  OA22X1_S38584 U6898 ( .IN1(g2436), .IN2(n1619), .IN3(n3543), .IN4(n3513), .Q(g27322) );
  OA22X1_S38584 U6899 ( .IN1(g2433), .IN2(n1618), .IN3(n3543), .IN4(n3523), .Q(g27308) );
  OA22X1_S38584 U6900 ( .IN1(g2444), .IN2(n1617), .IN3(n3543), .IN4(n3538), .Q(g27292) );
  OA22X1_S38584 U6901 ( .IN1(g1742), .IN2(n1616), .IN3(n3578), .IN4(n3530), .Q(g27302) );
  OA22X1_S38584 U6902 ( .IN1(g1739), .IN2(n1615), .IN3(n3578), .IN4(n3549), .Q(g27288) );
  OA22X1_S38584 U6903 ( .IN1(g1750), .IN2(n1614), .IN3(n3578), .IN4(n3573), .Q(g27275) );
  OA22X1_S38584 U6904 ( .IN1(g1048), .IN2(n1613), .IN3(n3614), .IN4(n3556), .Q(g27282) );
  OA22X1_S38584 U6905 ( .IN1(g1045), .IN2(n1612), .IN3(n3614), .IN4(n3584), .Q(g27271) );
  OA22X1_S38584 U6906 ( .IN1(g1056), .IN2(n1611), .IN3(n3614), .IN4(n3609), .Q(g27263) );
  OA22X1_S38584 U6907 ( .IN1(g361), .IN2(n1610), .IN3(n3648), .IN4(n3591), .Q(g27265)
         );
  OA22X1_S38584 U6908 ( .IN1(g358), .IN2(n1609), .IN3(n3648), .IN4(n3620), .Q(g27259)
         );
  OA22X1_S38584 U6909 ( .IN1(g369), .IN2(n1608), .IN3(n3648), .IN4(n3643), .Q(g27256)
         );
  OA22X1_S38584 U6910 ( .IN1(g2466), .IN2(n1619), .IN3(n3512), .IN4(n3513), .Q(g27342) );
  OA22X1_S38584 U6911 ( .IN1(g2463), .IN2(n1618), .IN3(n3512), .IN4(n3523), .Q(g27335) );
  OA22X1_S38584 U6912 ( .IN1(g2473), .IN2(n1617), .IN3(n3512), .IN4(n3538), .Q(g27324) );
  OA22X1_S38584 U6913 ( .IN1(g1772), .IN2(n1616), .IN3(n3529), .IN4(n3530), .Q(g27330) );
  OA22X1_S38584 U6914 ( .IN1(test_so58), .IN2(n1615), .IN3(n3529), .IN4(n3549), .Q(
        g27318) );
  OA22X1_S38584 U6915 ( .IN1(g1779), .IN2(n1614), .IN3(n3529), .IN4(n3573), .Q(g27304) );
  OA22X1_S38584 U6916 ( .IN1(g1078), .IN2(n1613), .IN3(n3555), .IN4(n3556), .Q(g27313) );
  OA22X1_S38584 U6917 ( .IN1(g1075), .IN2(n1612), .IN3(n3555), .IN4(n3584), .Q(g27298) );
  OA22X1_S38584 U6918 ( .IN1(g1085), .IN2(n1611), .IN3(n3555), .IN4(n3609), .Q(g27284) );
  OA22X1_S38584 U6919 ( .IN1(g391), .IN2(n1610), .IN3(n3590), .IN4(n3591), .Q(g27293)
         );
  OA22X1_S38584 U6920 ( .IN1(g388), .IN2(n1609), .IN3(n3590), .IN4(n3620), .Q(g27278)
         );
  OA22X1_S38584 U6921 ( .IN1(g398), .IN2(n1608), .IN3(n3590), .IN4(n3643), .Q(g27267)
         );
  OA22X1_S38584 U6922 ( .IN1(g2421), .IN2(n1619), .IN3(n3568), .IN4(n3513), .Q(g27307) );
  OA22X1_S38584 U6923 ( .IN1(g2418), .IN2(n1618), .IN3(n3568), .IN4(n3523), .Q(g27291) );
  OA22X1_S38584 U6924 ( .IN1(g2429), .IN2(n1617), .IN3(n3568), .IN4(n3538), .Q(g27276) );
  OA22X1_S38584 U6925 ( .IN1(g1727), .IN2(n1616), .IN3(n3604), .IN4(n3530), .Q(g27287) );
  OA22X1_S38584 U6926 ( .IN1(g1724), .IN2(n1615), .IN3(n3604), .IN4(n3549), .Q(g27274) );
  OA22X1_S38584 U6927 ( .IN1(g1735), .IN2(n1614), .IN3(n3604), .IN4(n3573), .Q(g27264) );
  OA22X1_S38584 U6928 ( .IN1(g1033), .IN2(n1613), .IN3(n3638), .IN4(n3556), .Q(g27270) );
  OA22X1_S38584 U6929 ( .IN1(g1030), .IN2(n1612), .IN3(n3638), .IN4(n3584), .Q(g27262) );
  OA22X1_S38584 U6930 ( .IN1(g1041), .IN2(n1611), .IN3(n3638), .IN4(n3609), .Q(g27257) );
  OA22X1_S38584 U6931 ( .IN1(test_so16), .IN2(n1610), .IN3(n3665), .IN4(n3591), .Q(
        g27258) );
  OA22X1_S38584 U6932 ( .IN1(g343), .IN2(n1609), .IN3(n3665), .IN4(n3620), .Q(g27255)
         );
  OA22X1_S38584 U6933 ( .IN1(g354), .IN2(n1608), .IN3(n3665), .IN4(n3643), .Q(g27253)
         );
  OA22X1_S38584 U6934 ( .IN1(n4731), .IN2(n4193), .IN3(g2878), .IN4(n4716), .Q(g21882) );
  NAND2X0 U6935 ( .IN1(n4194), .IN2(n4195), .QN(n4193) );
  OA22X1_S38584 U6936 ( .IN1(n4731), .IN2(n4196), .IN3(g2877), .IN4(n4716), .Q(g21880) );
  NAND2X0 U6937 ( .IN1(n4197), .IN2(n4198), .QN(n4196) );
  OA22X1_S38584 U6938 ( .IN1(g2479), .IN2(n3748), .IN3(n4664), .IN4(n3749), .Q(g26676) );
  NOR2X0 U6939 ( .IN1(n4524), .IN2(n4385), .QN(n3748) );
  OA22X1_S38584 U6940 ( .IN1(g2524), .IN2(n3438), .IN3(n4664), .IN4(n3436), .Q(g27769) );
  NOR2X0 U6941 ( .IN1(n3437), .IN2(n4524), .QN(n3438) );
  OA22X1_S38584 U6942 ( .IN1(g2503), .IN2(n3179), .IN3(n4664), .IN4(n3177), .Q(g28783) );
  NOR2X0 U6943 ( .IN1(n3178), .IN2(n4524), .QN(n3179) );
  OA22X1_S38584 U6944 ( .IN1(g1785), .IN2(n3756), .IN3(n4667), .IN4(n3751), .Q(g26670) );
  NOR2X0 U6945 ( .IN1(n4525), .IN2(n4386), .QN(n3756) );
  OA22X1_S38584 U6946 ( .IN1(g1830), .IN2(n3450), .IN3(n4667), .IN4(n3440), .Q(g27766) );
  NOR2X0 U6947 ( .IN1(n3441), .IN2(n4525), .QN(n3450) );
  OA22X1_S38584 U6948 ( .IN1(g1809), .IN2(n3187), .IN3(n4667), .IN4(n3182), .Q(g28772) );
  NOR2X0 U6949 ( .IN1(n3183), .IN2(n4525), .QN(n3187) );
  OA22X1_S38584 U6950 ( .IN1(g1091), .IN2(n3786), .IN3(n4672), .IN4(n3758), .Q(g26665) );
  NOR2X0 U6951 ( .IN1(n4671), .IN2(n4387), .QN(n3786) );
  OA22X1_S38584 U6952 ( .IN1(g1136), .IN2(n3462), .IN3(n4672), .IN4(n3452), .Q(g27763) );
  NOR2X0 U6953 ( .IN1(n3453), .IN2(n4671), .QN(n3462) );
  OA22X1_S38584 U6954 ( .IN1(g1115), .IN2(n3203), .IN3(n4672), .IN4(n3190), .Q(g28759) );
  NOR2X0 U6955 ( .IN1(n3191), .IN2(n4671), .QN(n3203) );
  OA22X1_S38584 U6956 ( .IN1(test_so82), .IN2(n3862), .IN3(n4663), .IN4(n3749), .Q(
        g26025) );
  NOR2X0 U6957 ( .IN1(n4509), .IN2(n4385), .QN(n3862) );
  OA22X1_S38584 U6958 ( .IN1(g2478), .IN2(n3752), .IN3(n4665), .IN4(n3749), .Q(g26672) );
  NOR2X0 U6959 ( .IN1(n4516), .IN2(n4385), .QN(n3752) );
  OA22X1_S38584 U6960 ( .IN1(test_so81), .IN2(n3435), .IN3(n4663), .IN4(n3436), .Q(
        g27771) );
  NOR2X0 U6961 ( .IN1(n3437), .IN2(n4509), .QN(n3435) );
  OA22X1_S38584 U6962 ( .IN1(g2523), .IN2(n3442), .IN3(n4665), .IN4(n3436), .Q(g27767) );
  NOR2X0 U6963 ( .IN1(n3437), .IN2(n4516), .QN(n3442) );
  OA22X1_S38584 U6964 ( .IN1(g2501), .IN2(n3176), .IN3(n4663), .IN4(n3177), .Q(g28788) );
  NOR2X0 U6965 ( .IN1(n3178), .IN2(n4509), .QN(n3176) );
  OA22X1_S38584 U6966 ( .IN1(g2502), .IN2(n3184), .IN3(n4665), .IN4(n3177), .Q(g28774) );
  NOR2X0 U6967 ( .IN1(n3178), .IN2(n4516), .QN(n3184) );
  OA22X1_S38584 U6968 ( .IN1(g1783), .IN2(n3750), .IN3(n4666), .IN4(n3751), .Q(g26675) );
  NOR2X0 U6969 ( .IN1(n4511), .IN2(n4386), .QN(n3750) );
  OA22X1_S38584 U6970 ( .IN1(test_so60), .IN2(n3759), .IN3(n4668), .IN4(n3751), .Q(
        g26667) );
  NOR2X0 U6971 ( .IN1(n4518), .IN2(n4386), .QN(n3759) );
  OA22X1_S38584 U6972 ( .IN1(g1828), .IN2(n3439), .IN3(n4666), .IN4(n3440), .Q(g27768) );
  NOR2X0 U6973 ( .IN1(n3441), .IN2(n4511), .QN(n3439) );
  OA22X1_S38584 U6974 ( .IN1(g1829), .IN2(n3454), .IN3(n4668), .IN4(n3440), .Q(g27764) );
  NOR2X0 U6975 ( .IN1(n3441), .IN2(n4518), .QN(n3454) );
  OA22X1_S38584 U6976 ( .IN1(g1807), .IN2(n3181), .IN3(n4666), .IN4(n3182), .Q(g28778) );
  NOR2X0 U6977 ( .IN1(n3183), .IN2(n4511), .QN(n3181) );
  OA22X1_S38584 U6978 ( .IN1(g1808), .IN2(n3200), .IN3(n4668), .IN4(n3182), .Q(g28761) );
  NOR2X0 U6979 ( .IN1(n3183), .IN2(n4518), .QN(n3200) );
  OA22X1_S38584 U6980 ( .IN1(g1089), .IN2(n3757), .IN3(n4670), .IN4(n3758), .Q(g26669) );
  NOR2X0 U6981 ( .IN1(n4669), .IN2(n4387), .QN(n3757) );
  OA22X1_S38584 U6982 ( .IN1(g1090), .IN2(n3789), .IN3(n4674), .IN4(n3758), .Q(g26661) );
  NOR2X0 U6983 ( .IN1(n4673), .IN2(n4387), .QN(n3789) );
  OA22X1_S38584 U6984 ( .IN1(g1134), .IN2(n3451), .IN3(n4670), .IN4(n3452), .Q(g27765) );
  NOR2X0 U6985 ( .IN1(n3453), .IN2(n4669), .QN(n3451) );
  OA22X1_S38584 U6986 ( .IN1(g1135), .IN2(n3466), .IN3(n4674), .IN4(n3452), .Q(g27761) );
  NOR2X0 U6987 ( .IN1(n3453), .IN2(n4673), .QN(n3466) );
  OA22X1_S38584 U6988 ( .IN1(g1113), .IN2(n3189), .IN3(n4670), .IN4(n3190), .Q(g28767) );
  NOR2X0 U6989 ( .IN1(n3191), .IN2(n4669), .QN(n3189) );
  OA22X1_S38584 U6990 ( .IN1(g1114), .IN2(n3216), .IN3(n4674), .IN4(n3190), .Q(g28747) );
  NOR2X0 U6991 ( .IN1(n3191), .IN2(n4673), .QN(n3216) );
  OA22X1_S38584 U6992 ( .IN1(g402), .IN2(n3787), .IN3(n4675), .IN4(n3788), .Q(g26664)
         );
  NOR2X0 U6993 ( .IN1(n4506), .IN2(n4388), .QN(n3787) );
  OA22X1_S38584 U6994 ( .IN1(g404), .IN2(n3816), .IN3(n4677), .IN4(n3788), .Q(g26659)
         );
  NOR2X0 U6995 ( .IN1(n4676), .IN2(n4388), .QN(n3816) );
  OA22X1_S38584 U6996 ( .IN1(g403), .IN2(n3817), .IN3(n4678), .IN4(n3788), .Q(g26655)
         );
  NOR2X0 U6997 ( .IN1(n4520), .IN2(n4388), .QN(n3817) );
  OA22X1_S38584 U6998 ( .IN1(g447), .IN2(n3463), .IN3(n4675), .IN4(n3464), .Q(g27762)
         );
  NOR2X0 U6999 ( .IN1(n3465), .IN2(n4506), .QN(n3463) );
  OA22X1_S38584 U7000 ( .IN1(g449), .IN2(n3474), .IN3(n4677), .IN4(n3464), .Q(g27760)
         );
  NOR2X0 U7001 ( .IN1(n3465), .IN2(n4676), .QN(n3474) );
  OA22X1_S38584 U7002 ( .IN1(g448), .IN2(n3475), .IN3(n4678), .IN4(n3464), .Q(g27759)
         );
  NOR2X0 U7003 ( .IN1(n3465), .IN2(n4520), .QN(n3475) );
  OA22X1_S38584 U7004 ( .IN1(g426), .IN2(n3205), .IN3(n4675), .IN4(n3206), .Q(g28754)
         );
  NOR2X0 U7005 ( .IN1(n3207), .IN2(n4506), .QN(n3205) );
  OA22X1_S38584 U7006 ( .IN1(g428), .IN2(n3219), .IN3(n4677), .IN4(n3206), .Q(g28745)
         );
  NOR2X0 U7007 ( .IN1(n3207), .IN2(n4676), .QN(n3219) );
  OA22X1_S38584 U7008 ( .IN1(test_so17), .IN2(n3230), .IN3(n4678), .IN4(n3206), .Q(
        g28736) );
  NOR2X0 U7009 ( .IN1(n3207), .IN2(n4520), .QN(n3230) );
  NBUFFX2 U7010 ( .IN(g2624), .Q(n4600) );
  NBUFFX2 U7011 ( .IN(g1930), .Q(n4612) );
  NBUFFX2 U7012 ( .IN(g1236), .Q(n4624) );
  NBUFFX2 U7013 ( .IN(g550), .Q(n4634) );
  OA21X1 U7014 ( .IN1(g2374), .IN2(DFF_1378_n1), .IN3(n2963), .Q(g30055) );
  AO221X1 U7015 ( .IN1(g28903), .IN2(n4608), .IN3(g2380), .IN4(n4524), .IN5(
        n4487), .Q(n2963) );
  NBUFFX2 U7016 ( .IN(g963), .Q(g5472) );
  NAND4X0 U7017 ( .IN1(g2165), .IN2(g2170), .IN3(n4035), .IN4(n4036), .QN(
        n3198) );
  NOR2X0 U7018 ( .IN1(n4389), .IN2(n4319), .QN(n4035) );
  NOR4X0 U7019 ( .IN1(n4287), .IN2(n4563), .IN3(n4555), .IN4(n4325), .QN(n4036) );
  NAND4X0 U7020 ( .IN1(g1471), .IN2(g1476), .IN3(n4041), .IN4(n4042), .QN(
        n3214) );
  NOR2X0 U7021 ( .IN1(n4390), .IN2(n4320), .QN(n4041) );
  NOR4X0 U7022 ( .IN1(n4288), .IN2(n4565), .IN3(n4557), .IN4(n4326), .QN(n4042) );
  NBUFFX2 U7023 ( .IN(g1088), .Q(n4630) );
  XOR2X1 U7024 ( .IN1(g8261), .IN2(g8260), .Q(n4230) );
  XOR2X1 U7025 ( .IN1(g8275), .IN2(g8274), .Q(n4226) );
  XOR2X1 U7026 ( .IN1(g2969), .IN2(test_so2), .Q(n4205) );
  XOR2X1 U7027 ( .IN1(g2944), .IN2(g2941), .Q(n4216) );
  XNOR2X1 U7028 ( .IN1(g2133), .IN2(n2501), .Q(n2493) );
  XNOR2X1 U7029 ( .IN1(g1439), .IN2(n2528), .Q(n2520) );
  XNOR2X1 U7030 ( .IN1(g753), .IN2(n2554), .Q(n2546) );
  XNOR2X1 U7031 ( .IN1(g65), .IN2(n2580), .Q(n2572) );
  XNOR2X1 U7032 ( .IN1(g2129), .IN2(n2502), .Q(n2492) );
  XNOR2X1 U7033 ( .IN1(g1435), .IN2(n2529), .Q(n2519) );
  XNOR2X1 U7034 ( .IN1(test_so36), .IN2(n2555), .Q(n2545) );
  XNOR2X1 U7035 ( .IN1(g61), .IN2(n2581), .Q(n2571) );
  XNOR2X1 U7036 ( .IN1(g2138), .IN2(n2503), .Q(n2491) );
  XNOR2X1 U7037 ( .IN1(g1444), .IN2(n2530), .Q(n2518) );
  XNOR2X1 U7038 ( .IN1(g758), .IN2(n2556), .Q(n2544) );
  XNOR2X1 U7039 ( .IN1(g70), .IN2(n2582), .Q(n2570) );
  NOR3X0 U7040 ( .IN1(n2508), .IN2(n2509), .IN3(n2510), .QN(n2507) );
  XOR2X1 U7041 ( .IN1(n2513), .IN2(g2160), .Q(n2508) );
  XNOR2X1 U7042 ( .IN1(n2511), .IN2(g2142), .Q(n2510) );
  XOR2X1 U7043 ( .IN1(n2512), .IN2(test_so78), .Q(n2509) );
  NOR3X0 U7044 ( .IN1(n2534), .IN2(n2535), .IN3(n2536), .QN(n2533) );
  XOR2X1 U7045 ( .IN1(n2539), .IN2(g1466), .Q(n2534) );
  XNOR2X1 U7046 ( .IN1(n2537), .IN2(g1448), .Q(n2536) );
  XOR2X1 U7047 ( .IN1(n2538), .IN2(g1462), .Q(n2535) );
  NOR3X0 U7048 ( .IN1(n2586), .IN2(n2587), .IN3(n2588), .QN(n2585) );
  XOR2X1 U7049 ( .IN1(n2591), .IN2(g92), .Q(n2586) );
  XNOR2X1 U7050 ( .IN1(n2589), .IN2(g74), .Q(n2588) );
  XOR2X1 U7051 ( .IN1(n2590), .IN2(g88), .Q(n2587) );
  NOR2X0 U7052 ( .IN1(n3704), .IN2(n3705), .QN(n3701) );
  NOR3X0 U7053 ( .IN1(n4405), .IN2(g185), .IN3(n3706), .QN(n3704) );
  NBUFFX2 U7054 ( .IN(g2987), .Q(n4595) );
  NOR3X0 U7055 ( .IN1(n2560), .IN2(n2561), .IN3(n2562), .QN(n2559) );
  XOR2X1 U7056 ( .IN1(n2565), .IN2(g780), .Q(n2560) );
  XNOR2X1 U7057 ( .IN1(n2563), .IN2(g762), .Q(n2562) );
  XOR2X1 U7058 ( .IN1(n2564), .IN2(g776), .Q(n2561) );
  NOR2X0 U7059 ( .IN1(n3969), .IN2(n3970), .QN(n3968) );
  XOR2X1 U7060 ( .IN1(n2154), .IN2(test_so92), .Q(n3969) );
  XOR2X1 U7061 ( .IN1(n2155), .IN2(g2753), .Q(n3970) );
  NOR2X0 U7062 ( .IN1(n3963), .IN2(n3964), .QN(n3962) );
  XOR2X1 U7063 ( .IN1(n2159), .IN2(g2707), .Q(n3963) );
  XOR2X1 U7064 ( .IN1(n2160), .IN2(g2727), .Q(n3964) );
  NOR2X0 U7065 ( .IN1(n3989), .IN2(n3990), .QN(n3988) );
  XOR2X1 U7066 ( .IN1(n2052), .IN2(g2046), .Q(n3989) );
  XOR2X1 U7067 ( .IN1(n2053), .IN2(g2059), .Q(n3990) );
  NOR2X0 U7068 ( .IN1(n3983), .IN2(n3984), .QN(n3982) );
  XOR2X1 U7069 ( .IN1(n2057), .IN2(g2013), .Q(n3983) );
  XOR2X1 U7070 ( .IN1(n2058), .IN2(g2033), .Q(n3984) );
  NOR2X0 U7071 ( .IN1(n4011), .IN2(n4012), .QN(n4010) );
  XOR2X1 U7072 ( .IN1(n1950), .IN2(g1352), .Q(n4011) );
  XOR2X1 U7073 ( .IN1(n1951), .IN2(g1365), .Q(n4012) );
  NOR2X0 U7074 ( .IN1(n4005), .IN2(n4006), .QN(n4004) );
  XOR2X1 U7075 ( .IN1(n1955), .IN2(g1319), .Q(n4005) );
  XOR2X1 U7076 ( .IN1(n1956), .IN2(g1339), .Q(n4006) );
  NOR2X0 U7077 ( .IN1(n4029), .IN2(n4030), .QN(n4028) );
  XOR2X1 U7078 ( .IN1(n1849), .IN2(test_so28), .Q(n4029) );
  XOR2X1 U7079 ( .IN1(n1850), .IN2(g679), .Q(n4030) );
  NOR2X0 U7080 ( .IN1(n4023), .IN2(n4024), .QN(n4022) );
  XOR2X1 U7081 ( .IN1(n1854), .IN2(g633), .Q(n4023) );
  XOR2X1 U7082 ( .IN1(n1855), .IN2(g653), .Q(n4024) );
  XOR2X1 U7083 ( .IN1(g2990), .IN2(n2420), .Q(N690) );
  XOR2X1 U7084 ( .IN1(g3083), .IN2(n2421), .Q(N995) );
  XOR2X1 U7085 ( .IN1(g2962), .IN2(n1629), .Q(n4281) );
  XOR2X1 U7086 ( .IN1(g2934), .IN2(n1628), .Q(n4280) );
  NOR2X0 U7087 ( .IN1(n2164), .IN2(n3413), .QN(g28328) );
  XOR2X1 U7088 ( .IN1(n3414), .IN2(g2766), .Q(n3413) );
  OR2X1 U7089 ( .IN1(n4393), .IN2(n3415), .Q(n3414) );
  NOR2X0 U7090 ( .IN1(n2164), .IN2(n3483), .QN(g27724) );
  XOR2X1 U7091 ( .IN1(n3415), .IN2(g2760), .Q(n3483) );
  NOR2X0 U7092 ( .IN1(n2164), .IN2(n3737), .QN(g26795) );
  XOR2X1 U7093 ( .IN1(n3681), .IN2(test_so92), .Q(n3737) );
  NOR2X0 U7094 ( .IN1(n2062), .IN2(n3416), .QN(g28325) );
  XOR2X1 U7095 ( .IN1(n3417), .IN2(g2072), .Q(n3416) );
  OR2X1 U7096 ( .IN1(n4394), .IN2(n3418), .Q(n3417) );
  NOR2X0 U7097 ( .IN1(n2062), .IN2(n3484), .QN(g27722) );
  XOR2X1 U7098 ( .IN1(n3418), .IN2(test_so70), .Q(n3484) );
  NOR2X0 U7099 ( .IN1(n2062), .IN2(n3738), .QN(g26789) );
  XOR2X1 U7100 ( .IN1(n3489), .IN2(g2046), .Q(n3738) );
  NOR2X0 U7101 ( .IN1(n1960), .IN2(n3419), .QN(g28321) );
  XOR2X1 U7102 ( .IN1(n3420), .IN2(g1378), .Q(n3419) );
  OR2X1 U7103 ( .IN1(n4395), .IN2(n3421), .Q(n3420) );
  NOR2X0 U7104 ( .IN1(n1960), .IN2(n3485), .QN(g27718) );
  XOR2X1 U7105 ( .IN1(n3421), .IN2(g1372), .Q(n3485) );
  NOR2X0 U7106 ( .IN1(n1960), .IN2(n3743), .QN(g26781) );
  XOR2X1 U7107 ( .IN1(n3493), .IN2(g1352), .Q(n3743) );
  NOR2X0 U7108 ( .IN1(n1859), .IN2(n3241), .QN(g28668) );
  XOR2X1 U7109 ( .IN1(n3242), .IN2(g692), .Q(n3241) );
  OR2X1 U7110 ( .IN1(n4396), .IN2(n3243), .Q(n3242) );
  NOR2X0 U7111 ( .IN1(n1859), .IN2(n3422), .QN(g28199) );
  XOR2X1 U7112 ( .IN1(n3243), .IN2(g686), .Q(n3422) );
  NOR2X0 U7113 ( .IN1(n1859), .IN2(n3744), .QN(g26776) );
  XOR2X1 U7114 ( .IN1(n3497), .IN2(test_so28), .Q(n3744) );
  NOR3X0 U7115 ( .IN1(n4057), .IN2(n3736), .IN3(n3734), .QN(g25201) );
  ISOLANDX1 U7116 ( .D(n4058), .ISO(g2903), .Q(n4057) );
  NOR3X0 U7117 ( .IN1(n4122), .IN2(n4059), .IN3(n3734), .QN(g23358) );
  ISOLANDX1 U7118 ( .D(n4123), .ISO(g2896), .Q(n4122) );
  NBUFFX2 U7119 ( .IN(g2950), .Q(n4649) );
  NOR2X0 U7120 ( .IN1(n1606), .IN2(n3244), .QN(g28637) );
  XOR2X1 U7121 ( .IN1(n3160), .IN2(g2133), .Q(n3244) );
  NOR2X0 U7122 ( .IN1(n1606), .IN2(n3498), .QN(g27621) );
  XOR2X1 U7123 ( .IN1(n4522), .IN2(g2142), .Q(n3498) );
  NOR2X0 U7124 ( .IN1(n1606), .IN2(n3850), .QN(g26532) );
  XOR2X1 U7125 ( .IN1(n4526), .IN2(g2151), .Q(n3850) );
  NOR2X0 U7126 ( .IN1(n1606), .IN2(n4069), .QN(g25067) );
  XOR2X1 U7127 ( .IN1(n3888), .IN2(g2160), .Q(n4069) );
  NOR2X0 U7128 ( .IN1(n1605), .IN2(n3245), .QN(g28636) );
  XOR2X1 U7129 ( .IN1(n3164), .IN2(g1439), .Q(n3245) );
  NOR2X0 U7130 ( .IN1(n1605), .IN2(n3499), .QN(g27612) );
  XOR2X1 U7131 ( .IN1(n4523), .IN2(g1448), .Q(n3499) );
  NOR2X0 U7132 ( .IN1(n1605), .IN2(n3851), .QN(g26531) );
  XOR2X1 U7133 ( .IN1(n4527), .IN2(g1457), .Q(n3851) );
  NOR2X0 U7134 ( .IN1(n1605), .IN2(n4070), .QN(g25056) );
  XOR2X1 U7135 ( .IN1(n3891), .IN2(g1466), .Q(n4070) );
  NOR2X0 U7136 ( .IN1(n1604), .IN2(n3246), .QN(g28635) );
  XOR2X1 U7137 ( .IN1(n3168), .IN2(g753), .Q(n3246) );
  NOR2X0 U7138 ( .IN1(n1604), .IN2(n3500), .QN(g27603) );
  XOR2X1 U7139 ( .IN1(n3431), .IN2(g762), .Q(n3500) );
  NOR2X0 U7140 ( .IN1(n1604), .IN2(n3852), .QN(g26530) );
  XOR2X1 U7141 ( .IN1(n3690), .IN2(g771), .Q(n3852) );
  NOR2X0 U7142 ( .IN1(n1604), .IN2(n4071), .QN(g25042) );
  XOR2X1 U7143 ( .IN1(n3894), .IN2(g780), .Q(n4071) );
  NOR2X0 U7144 ( .IN1(n1603), .IN2(n3247), .QN(g28634) );
  XOR2X1 U7145 ( .IN1(n3172), .IN2(g65), .Q(n3247) );
  NOR2X0 U7146 ( .IN1(n1603), .IN2(n3501), .QN(g27594) );
  XOR2X1 U7147 ( .IN1(n4521), .IN2(g74), .Q(n3501) );
  NOR2X0 U7148 ( .IN1(n1603), .IN2(n3853), .QN(g26529) );
  XOR2X1 U7149 ( .IN1(n4528), .IN2(g83), .Q(n3853) );
  NOR2X0 U7150 ( .IN1(n1603), .IN2(n4072), .QN(g25027) );
  XOR2X1 U7151 ( .IN1(n3897), .IN2(g92), .Q(n4072) );
  NOR2X0 U7152 ( .IN1(n1585), .IN2(n4060), .QN(g25199) );
  XOR2X1 U7153 ( .IN1(n4061), .IN2(g2920), .Q(n4060) );
  AOI21X1 U7154 ( .IN1(g1886), .IN2(DFF_1133_n1), .IN3(n3173), .QN(g28990) );
  OA221X1 U7155 ( .IN1(n4614), .IN2(DFF_1142_n1), .IN3(n4315), .IN4(n3174), 
        .IN5(n4493), .Q(n3173) );
  OA21X1 U7156 ( .IN1(n4581), .IN2(g1680), .IN3(n4582), .Q(g28903) );
  AO221X1 U7157 ( .IN1(n4525), .IN2(g1686), .IN3(n4620), .IN4(g26183), .IN5(
        n4488), .Q(n4582) );
  OA21X1 U7158 ( .IN1(n4583), .IN2(g986), .IN3(n4584), .Q(g26183) );
  AO221X1 U7159 ( .IN1(n4671), .IN2(g992), .IN3(g21346), .IN4(g6712), .IN5(
        n4432), .Q(n4584) );
  INVX0 U7160 ( .IN(g3234), .QN(n1582) );
  NAND2X0 U7161 ( .IN1(g7487), .IN2(n2148), .QN(n3951) );
  NAND2X0 U7162 ( .IN1(g7425), .IN2(n2148), .QN(n3954) );
  NAND2X0 U7163 ( .IN1(g7357), .IN2(n2046), .QN(n3971) );
  NAND2X0 U7164 ( .IN1(g7229), .IN2(n2046), .QN(n3974) );
  NAND2X0 U7165 ( .IN1(g7161), .IN2(n1944), .QN(n3991) );
  NAND2X0 U7166 ( .IN1(g6979), .IN2(n1944), .QN(n3996) );
  NAND2X0 U7167 ( .IN1(g6911), .IN2(n1843), .QN(n4013) );
  NAND2X0 U7168 ( .IN1(g6677), .IN2(n1843), .QN(n4014) );
  NAND2X0 U7169 ( .IN1(g2703), .IN2(n2148), .QN(n3950) );
  NAND2X0 U7170 ( .IN1(g2009), .IN2(n2046), .QN(n3953) );
  NAND2X0 U7171 ( .IN1(g1315), .IN2(n1944), .QN(n3973) );
  NAND2X0 U7172 ( .IN1(g629), .IN2(n1843), .QN(n3993) );
  NAND2X0 U7173 ( .IN1(g2704), .IN2(g7487), .QN(n3678) );
  NAND2X0 U7174 ( .IN1(g2010), .IN2(g7357), .QN(n3486) );
  NAND2X0 U7175 ( .IN1(g1316), .IN2(g7161), .QN(n3490) );
  NAND2X0 U7176 ( .IN1(g630), .IN2(g6911), .QN(n3494) );
  NAND2X0 U7177 ( .IN1(g2257), .IN2(g7084), .QN(n4170) );
  NAND2X0 U7178 ( .IN1(g2257), .IN2(g2214), .QN(n4172) );
  NAND2X0 U7179 ( .IN1(g1563), .IN2(n4589), .QN(n4173) );
  NAND2X0 U7180 ( .IN1(g1563), .IN2(g1520), .QN(n4175) );
  NAND2X0 U7181 ( .IN1(g869), .IN2(n4591), .QN(n4176) );
  NAND2X0 U7182 ( .IN1(g869), .IN2(n4592), .QN(n4178) );
  NAND2X0 U7183 ( .IN1(g181), .IN2(g6313), .QN(n4179) );
  NAND2X0 U7184 ( .IN1(g181), .IN2(g138), .QN(n4180) );
  NAND2X0 U7185 ( .IN1(g2704), .IN2(g7425), .QN(n4153) );
  NAND2X0 U7186 ( .IN1(g2010), .IN2(g7229), .QN(n4159) );
  NAND2X0 U7187 ( .IN1(g1316), .IN2(g6979), .QN(n4165) );
  NAND2X0 U7188 ( .IN1(g630), .IN2(g6677), .QN(n4168) );
  NOR2X0 U7189 ( .IN1(n4425), .IN2(g3231), .QN(n4200) );
  NAND2X0 U7190 ( .IN1(g2704), .IN2(g2703), .QN(n4146) );
  NAND2X0 U7191 ( .IN1(g2010), .IN2(g2009), .QN(n4150) );
  NAND2X0 U7192 ( .IN1(g1316), .IN2(g1315), .QN(n4156) );
  NAND2X0 U7193 ( .IN1(g630), .IN2(g629), .QN(n4162) );
  NAND3X0 U7194 ( .IN1(g2599), .IN2(n4426), .IN3(g2612), .QN(n4147) );
  NAND3X0 U7195 ( .IN1(g1905), .IN2(n4427), .IN3(test_so69), .QN(n4151) );
  NAND3X0 U7196 ( .IN1(g1211), .IN2(n4428), .IN3(g1224), .QN(n4157) );
  NAND3X0 U7197 ( .IN1(g525), .IN2(n4429), .IN3(g538), .QN(n4163) );
  NOR4X0 U7198 ( .IN1(n4327), .IN2(n4289), .IN3(g805), .IN4(g809), .QN(n4050)
         );
  NOR4X0 U7199 ( .IN1(n4328), .IN2(n4290), .IN3(g117), .IN4(g121), .QN(n4054)
         );
  NOR4X0 U7200 ( .IN1(n4325), .IN2(n4287), .IN3(g2190), .IN4(g2195), .QN(n4039) );
  NOR4X0 U7201 ( .IN1(n4326), .IN2(n4288), .IN3(g1496), .IN4(g1501), .QN(n4045) );
  OA222X1 U7202 ( .IN1(g2562), .IN2(n4299), .IN3(test_so87), .IN4(n4314), 
        .IN5(g2561), .IN6(n4370), .Q(g13194) );
  OA222X1 U7203 ( .IN1(g2559), .IN2(n4299), .IN3(g2539), .IN4(n4314), .IN5(
        g2555), .IN6(n4370), .Q(g13143) );
  OA222X1 U7204 ( .IN1(g2553), .IN2(n4299), .IN3(g2554), .IN4(n4314), .IN5(
        g2552), .IN6(n4370), .Q(g13175) );
  OA222X1 U7205 ( .IN1(g1868), .IN2(n4366), .IN3(g1869), .IN4(n4296), .IN5(
        g1867), .IN6(n4315), .Q(g13182) );
  OA222X1 U7206 ( .IN1(g1865), .IN2(n4366), .IN3(g1845), .IN4(n4296), .IN5(
        g1861), .IN6(n4315), .Q(g13135) );
  OA222X1 U7207 ( .IN1(g1859), .IN2(n4366), .IN3(g1860), .IN4(n4296), .IN5(
        g1858), .IN6(n4315), .Q(g13164) );
  OA222X1 U7208 ( .IN1(test_so44), .IN2(n4300), .IN3(g1175), .IN4(n4371), 
        .IN5(g1173), .IN6(n4316), .Q(g13171) );
  OA222X1 U7209 ( .IN1(g1171), .IN2(n4300), .IN3(g1151), .IN4(n4371), .IN5(
        g1167), .IN6(n4316), .Q(g13124) );
  OA222X1 U7210 ( .IN1(g1165), .IN2(n4300), .IN3(g1166), .IN4(n4371), .IN5(
        g1164), .IN6(n4316), .Q(g13155) );
  OA222X1 U7211 ( .IN1(g487), .IN2(n4313), .IN3(g488), .IN4(n4298), .IN5(g486), 
        .IN6(n4372), .Q(g13160) );
  OA222X1 U7212 ( .IN1(g484), .IN2(n4313), .IN3(g464), .IN4(n4298), .IN5(g480), 
        .IN6(n4372), .Q(g13111) );
  OA222X1 U7213 ( .IN1(g478), .IN2(n4313), .IN3(g479), .IN4(n4298), .IN5(g477), 
        .IN6(n4372), .Q(g13149) );
  AND3X1 U7214 ( .IN1(n3747), .IN2(n3678), .IN3(n4104), .Q(g24438) );
  OR2X1 U7215 ( .IN1(n4105), .IN2(g2720), .Q(n4104) );
  AND3X1 U7216 ( .IN1(n3755), .IN2(n3486), .IN3(n4107), .Q(g24434) );
  OR2X1 U7217 ( .IN1(n4108), .IN2(g2026), .Q(n4107) );
  AND3X1 U7218 ( .IN1(n3785), .IN2(n3490), .IN3(n4110), .Q(g24430) );
  OR2X1 U7219 ( .IN1(n4111), .IN2(g1332), .Q(n4110) );
  AND3X1 U7220 ( .IN1(n3815), .IN2(n3494), .IN3(n4113), .Q(g24426) );
  OR2X1 U7221 ( .IN1(n4114), .IN2(g646), .Q(n4113) );
  AND3X1 U7222 ( .IN1(n4106), .IN2(n3678), .IN3(n4184), .Q(g21974) );
  OR2X1 U7223 ( .IN1(n4185), .IN2(g2707), .Q(n4184) );
  AND3X1 U7224 ( .IN1(n4109), .IN2(n3486), .IN3(n4187), .Q(g21972) );
  OR2X1 U7225 ( .IN1(n4188), .IN2(g2013), .Q(n4187) );
  AND3X1 U7226 ( .IN1(n4112), .IN2(n3490), .IN3(n4190), .Q(g21969) );
  OR2X1 U7227 ( .IN1(n4191), .IN2(g1319), .Q(n4190) );
  AND3X1 U7228 ( .IN1(n4115), .IN2(n3494), .IN3(n4133), .Q(g23136) );
  OR2X1 U7229 ( .IN1(n4134), .IN2(g633), .Q(n4133) );
  AO22X1 U7230 ( .IN1(test_so8), .IN2(n4494), .IN3(n4644), .IN4(g1880), .Q(
        g17383) );
  AO22X1 U7231 ( .IN1(g3176), .IN2(n4383), .IN3(n4646), .IN4(g1880), .Q(g17303) );
  AO22X1 U7232 ( .IN1(g3173), .IN2(n4382), .IN3(g8106), .IN4(g1880), .Q(g17248) );
  AO22X1 U7233 ( .IN1(g3088), .IN2(n4494), .IN3(n4644), .IN4(g2574), .Q(g17429) );
  AO22X1 U7234 ( .IN1(g3185), .IN2(n4383), .IN3(n4646), .IN4(g2574), .Q(g17341) );
  AO22X1 U7235 ( .IN1(g3182), .IN2(n4382), .IN3(n4648), .IN4(g2574), .Q(g17271) );
  AO22X1 U7236 ( .IN1(n4644), .IN2(g499), .IN3(g3161), .IN4(n4494), .Q(g17302)
         );
  AO22X1 U7237 ( .IN1(n4646), .IN2(g499), .IN3(g3158), .IN4(n4383), .Q(g17247)
         );
  AO22X1 U7238 ( .IN1(n4648), .IN2(g499), .IN3(g3155), .IN4(n4382), .Q(g17229)
         );
  AO22X1 U7239 ( .IN1(n4600), .IN2(g2631), .IN3(g2584), .IN4(n4299), .Q(g18820) );
  AO22X1 U7240 ( .IN1(n4612), .IN2(g1937), .IN3(g1890), .IN4(n4366), .Q(g18794) );
  AO22X1 U7241 ( .IN1(n4624), .IN2(g1243), .IN3(g1196), .IN4(n4300), .Q(g18763) );
  AO22X1 U7242 ( .IN1(n4634), .IN2(g557), .IN3(test_so22), .IN4(n4313), .Q(
        g18726) );
  AO22X1 U7243 ( .IN1(g559), .IN2(g8106), .IN3(test_so6), .IN4(n4382), .Q(
        g18669) );
  AO22X1 U7244 ( .IN1(g559), .IN2(n4644), .IN3(g3084), .IN4(n4494), .Q(g18782)
         );
  AO22X1 U7245 ( .IN1(g559), .IN2(n4646), .IN3(g3211), .IN4(n4383), .Q(g18719)
         );
  AO22X1 U7246 ( .IN1(g2704), .IN2(n4292), .IN3(g2703), .IN4(g2584), .Q(g16718) );
  AO22X1 U7247 ( .IN1(g2010), .IN2(n4293), .IN3(g2009), .IN4(g1890), .Q(g16692) );
  AO22X1 U7248 ( .IN1(g1316), .IN2(n4294), .IN3(g1315), .IN4(g1196), .Q(g16671) );
  AO22X1 U7249 ( .IN1(g630), .IN2(n4295), .IN3(g629), .IN4(test_so22), .Q(
        g16654) );
  AO22X1 U7250 ( .IN1(g3170), .IN2(n4494), .IN3(n4644), .IN4(g1186), .Q(g17340) );
  AO22X1 U7251 ( .IN1(g3167), .IN2(n4383), .IN3(n4646), .IN4(g1186), .Q(g17270) );
  AO22X1 U7252 ( .IN1(g3164), .IN2(n4382), .IN3(n4648), .IN4(g1186), .Q(g17236) );
  AO22X1 U7253 ( .IN1(g2997), .IN2(n4596), .IN3(g3061), .IN4(n4365), .Q(g18907) );
  AO22X1 U7254 ( .IN1(g3078), .IN2(n4596), .IN3(g3060), .IN4(n4365), .Q(g18868) );
  AO22X1 U7255 ( .IN1(g3077), .IN2(n4596), .IN3(g3059), .IN4(n4365), .Q(g18837) );
  AO22X1 U7256 ( .IN1(g3076), .IN2(n4596), .IN3(g3058), .IN4(n4365), .Q(g18804) );
  AO22X1 U7257 ( .IN1(g3075), .IN2(n4596), .IN3(g3057), .IN4(n4365), .Q(g18755) );
  AO22X1 U7258 ( .IN1(g3074), .IN2(n4596), .IN3(g3056), .IN4(n4365), .Q(g16880) );
  AO22X1 U7259 ( .IN1(g3073), .IN2(n4596), .IN3(test_so96), .IN4(n4365), .Q(
        g16861) );
  AO22X1 U7260 ( .IN1(g3072), .IN2(n4596), .IN3(g3053), .IN4(n4365), .Q(g16854) );
  AO22X1 U7261 ( .IN1(g3071), .IN2(n4596), .IN3(g3052), .IN4(n4365), .Q(g16845) );
  AO22X1 U7262 ( .IN1(test_so97), .IN2(n4596), .IN3(g3051), .IN4(n4365), .Q(
        g16866) );
  AO22X1 U7263 ( .IN1(g3069), .IN2(n4596), .IN3(g3050), .IN4(n4365), .Q(g16857) );
  AO22X1 U7264 ( .IN1(g3068), .IN2(n4596), .IN3(g3049), .IN4(n4365), .Q(g16851) );
  AO22X1 U7265 ( .IN1(g3065), .IN2(n4596), .IN3(g3046), .IN4(n4365), .Q(g16860) );
  AO22X1 U7266 ( .IN1(g3064), .IN2(n4596), .IN3(g3045), .IN4(n4365), .Q(g16853) );
  AO22X1 U7267 ( .IN1(g3063), .IN2(n4596), .IN3(g3044), .IN4(n4365), .Q(g16844) );
  AO22X1 U7268 ( .IN1(g3091), .IN2(n4382), .IN3(g1939), .IN4(n4648), .Q(g17224) );
  AO22X1 U7269 ( .IN1(g3096), .IN2(n4494), .IN3(g2633), .IN4(n4644), .Q(g17269) );
  AO22X1 U7270 ( .IN1(g3093), .IN2(n4494), .IN3(g1939), .IN4(n4644), .Q(g17246) );
  AO22X1 U7271 ( .IN1(g3087), .IN2(n4494), .IN3(g1245), .IN4(n4644), .Q(g17234) );
  AO22X1 U7272 ( .IN1(g3067), .IN2(n4595), .IN3(g3048), .IN4(n4365), .Q(g16835) );
  AO22X1 U7273 ( .IN1(g3066), .IN2(n4595), .IN3(g3047), .IN4(n4365), .Q(g16803) );
  AO22X1 U7274 ( .IN1(g3062), .IN2(n4595), .IN3(g3043), .IN4(n4365), .Q(g16824) );
  AO22X1 U7275 ( .IN1(g3095), .IN2(n4383), .IN3(g2633), .IN4(n4646), .Q(g17235) );
  AO22X1 U7276 ( .IN1(g3094), .IN2(n4382), .IN3(g2633), .IN4(g8106), .Q(g17226) );
  AO22X1 U7277 ( .IN1(g3092), .IN2(n4383), .IN3(g1939), .IN4(n4646), .Q(g17228) );
  AO22X1 U7278 ( .IN1(g3086), .IN2(n4383), .IN3(g1245), .IN4(n4646), .Q(g17225) );
  AO22X1 U7279 ( .IN1(g3085), .IN2(n4382), .IN3(g1245), .IN4(g8106), .Q(g17222) );
  AO22X1 U7280 ( .IN1(g3099), .IN2(n4494), .IN3(n4644), .IN4(g21851), .Q(
        g25452) );
  AO22X1 U7281 ( .IN1(g3098), .IN2(n4383), .IN3(n4646), .IN4(g21851), .Q(
        g25451) );
  AO22X1 U7282 ( .IN1(g3097), .IN2(n4382), .IN3(g8106), .IN4(g21851), .Q(
        g25450) );
  NOR2X0 U7283 ( .IN1(n4586), .IN2(DFF_1_n1), .QN(g16823) );
  NOR2X0 U7284 ( .IN1(n3733), .IN2(n3734), .QN(g26798) );
  XOR2X1 U7285 ( .IN1(n3735), .IN2(g2908), .Q(n3733) );
  NAND2X0 U7286 ( .IN1(g2900), .IN2(n3736), .QN(n3735) );
  NOR2X0 U7287 ( .IN1(n4100), .IN2(n3734), .QN(g24473) );
  XNOR2X1 U7288 ( .IN1(n4059), .IN2(g2892), .Q(n4100) );
  NOR2X0 U7289 ( .IN1(n4181), .IN2(n3734), .QN(g22026) );
  XNOR2X1 U7290 ( .IN1(n2486), .IN2(g2888), .Q(n4181) );
  NAND2X0 U7291 ( .IN1(n4059), .IN2(g2892), .QN(n4058) );
  NAND2X0 U7292 ( .IN1(n2486), .IN2(g2888), .QN(n4123) );
  ISOLANDX1 U7293 ( .D(n4597), .ISO(g3234), .Q(g20877) );
  OA22X1_S38584 U7294 ( .IN1(g2801), .IN2(n2146), .IN3(n4415), .IN4(n3951), .Q(g20941) );
  OA22X1_S38584 U7295 ( .IN1(g2800), .IN2(n2145), .IN3(n4415), .IN4(n3954), .Q(g20919) );
  OA22X1_S38584 U7296 ( .IN1(g2798), .IN2(n2146), .IN3(n4393), .IN4(n3951), .Q(g21082) );
  OA22X1_S38584 U7297 ( .IN1(g2797), .IN2(n2145), .IN3(n4393), .IN4(n3954), .Q(g21075) );
  OA22X1_S38584 U7298 ( .IN1(g2795), .IN2(n2146), .IN3(n4471), .IN4(n3951), .Q(g21074) );
  OA22X1_S38584 U7299 ( .IN1(g2794), .IN2(n2145), .IN3(n4471), .IN4(n3954), .Q(g21062) );
  OA22X1_S38584 U7300 ( .IN1(g2792), .IN2(n2146), .IN3(n4467), .IN4(n3951), .Q(g21061) );
  OA22X1_S38584 U7301 ( .IN1(g2791), .IN2(n2145), .IN3(n4467), .IN4(n3954), .Q(g21045) );
  OA22X1_S38584 U7302 ( .IN1(g2789), .IN2(n2146), .IN3(n4407), .IN4(n3951), .Q(g21044) );
  OA22X1_S38584 U7303 ( .IN1(g2788), .IN2(n2145), .IN3(n4407), .IN4(n3954), .Q(g21027) );
  OA22X1_S38584 U7304 ( .IN1(g2786), .IN2(n2146), .IN3(n4397), .IN4(n3951), .Q(g21026) );
  OA22X1_S38584 U7305 ( .IN1(g2785), .IN2(n2145), .IN3(n4397), .IN4(n3954), .Q(g21006) );
  OA22X1_S38584 U7306 ( .IN1(g2783), .IN2(n2146), .IN3(n4408), .IN4(n3951), .Q(g21005) );
  OA22X1_S38584 U7307 ( .IN1(g2782), .IN2(n2145), .IN3(n4408), .IN4(n3954), .Q(g20983) );
  OA22X1_S38584 U7308 ( .IN1(g2780), .IN2(n2146), .IN3(n4419), .IN4(n3951), .Q(g20982) );
  OA22X1_S38584 U7309 ( .IN1(g2779), .IN2(n2145), .IN3(n4419), .IN4(n3954), .Q(g20964) );
  OA22X1_S38584 U7310 ( .IN1(g2777), .IN2(n2146), .IN3(n4472), .IN4(n3951), .Q(g20963) );
  OA22X1_S38584 U7311 ( .IN1(g2776), .IN2(n2145), .IN3(n4472), .IN4(n3954), .Q(g20940) );
  OA22X1_S38584 U7312 ( .IN1(g2774), .IN2(n2146), .IN3(n4398), .IN4(n3951), .Q(g20939) );
  OA22X1_S38584 U7313 ( .IN1(g2773), .IN2(n2145), .IN3(n4398), .IN4(n3954), .Q(g20918) );
  OA22X1_S38584 U7314 ( .IN1(test_so72), .IN2(n2044), .IN3(n4416), .IN4(n3971), .Q(
        g20917) );
  OA22X1_S38584 U7315 ( .IN1(g2106), .IN2(n2043), .IN3(n4416), .IN4(n3974), .Q(g20900) );
  OA22X1_S38584 U7316 ( .IN1(g2104), .IN2(n2044), .IN3(n4394), .IN4(n3971), .Q(g21072) );
  OA22X1_S38584 U7317 ( .IN1(g2103), .IN2(n2043), .IN3(n4394), .IN4(n3974), .Q(g21056) );
  OA22X1_S38584 U7318 ( .IN1(g2101), .IN2(n2044), .IN3(n4473), .IN4(n3971), .Q(g21055) );
  OA22X1_S38584 U7319 ( .IN1(g2100), .IN2(n2043), .IN3(n4473), .IN4(n3974), .Q(g21041) );
  OA22X1_S38584 U7320 ( .IN1(g2098), .IN2(n2044), .IN3(n4468), .IN4(n3971), .Q(g21040) );
  OA22X1_S38584 U7321 ( .IN1(g2097), .IN2(n2043), .IN3(n4468), .IN4(n3974), .Q(g21021) );
  OA22X1_S38584 U7322 ( .IN1(g2095), .IN2(n2044), .IN3(n4409), .IN4(n3971), .Q(g21020) );
  OA22X1_S38584 U7323 ( .IN1(g2094), .IN2(n2043), .IN3(n4409), .IN4(n3974), .Q(g21001) );
  OA22X1_S38584 U7324 ( .IN1(test_so71), .IN2(n2044), .IN3(n4399), .IN4(n3971), .Q(
        g21000) );
  OA22X1_S38584 U7325 ( .IN1(g2091), .IN2(n2043), .IN3(n4399), .IN4(n3974), .Q(g20979) );
  OA22X1_S38584 U7326 ( .IN1(g2089), .IN2(n2044), .IN3(n4410), .IN4(n3971), .Q(g20978) );
  OA22X1_S38584 U7327 ( .IN1(g2088), .IN2(n2043), .IN3(n4410), .IN4(n3974), .Q(g20955) );
  OA22X1_S38584 U7328 ( .IN1(g2086), .IN2(n2044), .IN3(n4420), .IN4(n3971), .Q(g20954) );
  OA22X1_S38584 U7329 ( .IN1(g2085), .IN2(n2043), .IN3(n4420), .IN4(n3974), .Q(g20936) );
  OA22X1_S38584 U7330 ( .IN1(g2083), .IN2(n2044), .IN3(n4474), .IN4(n3971), .Q(g20935) );
  OA22X1_S38584 U7331 ( .IN1(g2082), .IN2(n2043), .IN3(n4474), .IN4(n3974), .Q(g20916) );
  OA22X1_S38584 U7332 ( .IN1(g2080), .IN2(n2044), .IN3(n4400), .IN4(n3971), .Q(g20915) );
  OA22X1_S38584 U7333 ( .IN1(g2079), .IN2(n2043), .IN3(n4400), .IN4(n3974), .Q(g20899) );
  OA22X1_S38584 U7334 ( .IN1(g1413), .IN2(n1942), .IN3(n4417), .IN4(n3991), .Q(g20898) );
  OA22X1_S38584 U7335 ( .IN1(g1412), .IN2(n1941), .IN3(n4417), .IN4(n3996), .Q(g20883) );
  OA22X1_S38584 U7336 ( .IN1(g1410), .IN2(n1942), .IN3(n4395), .IN4(n3991), .Q(g21053) );
  OA22X1_S38584 U7337 ( .IN1(g1409), .IN2(n1941), .IN3(n4395), .IN4(n3996), .Q(g21035) );
  OA22X1_S38584 U7338 ( .IN1(g1407), .IN2(n1942), .IN3(n4475), .IN4(n3991), .Q(g21034) );
  OA22X1_S38584 U7339 ( .IN1(g1406), .IN2(n1941), .IN3(n4475), .IN4(n3996), .Q(g21017) );
  OA22X1_S38584 U7340 ( .IN1(g1404), .IN2(n1942), .IN3(n4469), .IN4(n3991), .Q(g21016) );
  OA22X1_S38584 U7341 ( .IN1(g1403), .IN2(n1941), .IN3(n4469), .IN4(n3996), .Q(g20995) );
  OA22X1_S38584 U7342 ( .IN1(test_so50), .IN2(n1942), .IN3(n4411), .IN4(n3991), .Q(
        g20994) );
  OA22X1_S38584 U7343 ( .IN1(g1400), .IN2(n1941), .IN3(n4411), .IN4(n3996), .Q(g20974) );
  OA22X1_S38584 U7344 ( .IN1(g1398), .IN2(n1942), .IN3(n4401), .IN4(n3991), .Q(g20973) );
  OA22X1_S38584 U7345 ( .IN1(g1397), .IN2(n1941), .IN3(n4401), .IN4(n3996), .Q(g20951) );
  OA22X1_S38584 U7346 ( .IN1(g1395), .IN2(n1942), .IN3(n4412), .IN4(n3991), .Q(g20950) );
  OA22X1_S38584 U7347 ( .IN1(g1394), .IN2(n1941), .IN3(n4412), .IN4(n3996), .Q(g20927) );
  OA22X1_S38584 U7348 ( .IN1(g1392), .IN2(n1942), .IN3(n4421), .IN4(n3991), .Q(g20926) );
  OA22X1_S38584 U7349 ( .IN1(g1391), .IN2(n1941), .IN3(n4421), .IN4(n3996), .Q(g20912) );
  OA22X1_S38584 U7350 ( .IN1(g1389), .IN2(n1942), .IN3(n4476), .IN4(n3991), .Q(g20911) );
  OA22X1_S38584 U7351 ( .IN1(g1388), .IN2(n1941), .IN3(n4476), .IN4(n3996), .Q(g20897) );
  OA22X1_S38584 U7352 ( .IN1(g1386), .IN2(n1942), .IN3(n4402), .IN4(n3991), .Q(g20896) );
  OA22X1_S38584 U7353 ( .IN1(test_so49), .IN2(n1941), .IN3(n4402), .IN4(n3996), .Q(
        g20882) );
  OA22X1_S38584 U7354 ( .IN1(test_so30), .IN2(n1841), .IN3(n4418), .IN4(n4013), .Q(
        g20881) );
  OA22X1_S38584 U7355 ( .IN1(g726), .IN2(n1840), .IN3(n4418), .IN4(n4014), .Q(g20876)
         );
  OA22X1_S38584 U7356 ( .IN1(g724), .IN2(n1841), .IN3(n4396), .IN4(n4013), .Q(g21032)
         );
  OA22X1_S38584 U7357 ( .IN1(g723), .IN2(n1840), .IN3(n4396), .IN4(n4014), .Q(g21011)
         );
  OA22X1_S38584 U7358 ( .IN1(g721), .IN2(n1841), .IN3(n4477), .IN4(n4013), .Q(g21010)
         );
  OA22X1_S38584 U7359 ( .IN1(g720), .IN2(n1840), .IN3(n4477), .IN4(n4014), .Q(g20991)
         );
  OA22X1_S38584 U7360 ( .IN1(g718), .IN2(n1841), .IN3(n4470), .IN4(n4013), .Q(g20990)
         );
  OA22X1_S38584 U7361 ( .IN1(g717), .IN2(n1840), .IN3(n4470), .IN4(n4014), .Q(g20968)
         );
  OA22X1_S38584 U7362 ( .IN1(g715), .IN2(n1841), .IN3(n4413), .IN4(n4013), .Q(g20967)
         );
  OA22X1_S38584 U7363 ( .IN1(g714), .IN2(n1840), .IN3(n4413), .IN4(n4014), .Q(g20946)
         );
  OA22X1_S38584 U7364 ( .IN1(g712), .IN2(n1841), .IN3(n4403), .IN4(n4013), .Q(g20945)
         );
  OA22X1_S38584 U7365 ( .IN1(test_so29), .IN2(n1840), .IN3(n4403), .IN4(n4014), .Q(
        g20923) );
  OA22X1_S38584 U7366 ( .IN1(g709), .IN2(n1841), .IN3(n4414), .IN4(n4013), .Q(g20922)
         );
  OA22X1_S38584 U7367 ( .IN1(g708), .IN2(n1840), .IN3(n4414), .IN4(n4014), .Q(g20903)
         );
  OA22X1_S38584 U7368 ( .IN1(g706), .IN2(n1841), .IN3(n4422), .IN4(n4013), .Q(g20902)
         );
  OA22X1_S38584 U7369 ( .IN1(g705), .IN2(n1840), .IN3(n4422), .IN4(n4014), .Q(g20893)
         );
  OA22X1_S38584 U7370 ( .IN1(g703), .IN2(n1841), .IN3(n4478), .IN4(n4013), .Q(g20892)
         );
  OA22X1_S38584 U7371 ( .IN1(g702), .IN2(n1840), .IN3(n4478), .IN4(n4014), .Q(g20880)
         );
  OA22X1_S38584 U7372 ( .IN1(g700), .IN2(n1841), .IN3(n4404), .IN4(n4013), .Q(g20879)
         );
  OA22X1_S38584 U7373 ( .IN1(g699), .IN2(n1840), .IN3(n4404), .IN4(n4014), .Q(g20875)
         );
  OA22X1_S38584 U7374 ( .IN1(g2799), .IN2(n2147), .IN3(n4415), .IN4(n3950), .Q(g20965) );
  OA22X1_S38584 U7375 ( .IN1(test_so94), .IN2(n2147), .IN3(n4393), .IN4(n3950), .Q(
        g21094) );
  OA22X1_S38584 U7376 ( .IN1(g2793), .IN2(n2147), .IN3(n4471), .IN4(n3950), .Q(g21081) );
  OA22X1_S38584 U7377 ( .IN1(g2790), .IN2(n2147), .IN3(n4467), .IN4(n3950), .Q(g21073) );
  OA22X1_S38584 U7378 ( .IN1(g2787), .IN2(n2147), .IN3(n4407), .IN4(n3950), .Q(g21060) );
  OA22X1_S38584 U7379 ( .IN1(g2784), .IN2(n2147), .IN3(n4397), .IN4(n3950), .Q(g21043) );
  OA22X1_S38584 U7380 ( .IN1(test_so93), .IN2(n2147), .IN3(n4408), .IN4(n3950), .Q(
        g21025) );
  OA22X1_S38584 U7381 ( .IN1(g2778), .IN2(n2147), .IN3(n4419), .IN4(n3950), .Q(g21004) );
  OA22X1_S38584 U7382 ( .IN1(g2775), .IN2(n2147), .IN3(n4472), .IN4(n3950), .Q(g20981) );
  OA22X1_S38584 U7383 ( .IN1(g2772), .IN2(n2147), .IN3(n4398), .IN4(n3950), .Q(g20962) );
  OA22X1_S38584 U7384 ( .IN1(g2105), .IN2(n2045), .IN3(n4416), .IN4(n3953), .Q(g20937) );
  OA22X1_S38584 U7385 ( .IN1(g2102), .IN2(n2045), .IN3(n4394), .IN4(n3953), .Q(g21080) );
  OA22X1_S38584 U7386 ( .IN1(g2099), .IN2(n2045), .IN3(n4473), .IN4(n3953), .Q(g21071) );
  OA22X1_S38584 U7387 ( .IN1(g2096), .IN2(n2045), .IN3(n4468), .IN4(n3953), .Q(g21054) );
  OA22X1_S38584 U7388 ( .IN1(g2093), .IN2(n2045), .IN3(n4409), .IN4(n3953), .Q(g21039) );
  OA22X1_S38584 U7389 ( .IN1(g2090), .IN2(n2045), .IN3(n4399), .IN4(n3953), .Q(g21019) );
  OA22X1_S38584 U7390 ( .IN1(g2087), .IN2(n2045), .IN3(n4410), .IN4(n3953), .Q(g20999) );
  OA22X1_S38584 U7391 ( .IN1(g2084), .IN2(n2045), .IN3(n4420), .IN4(n3953), .Q(g20977) );
  OA22X1_S38584 U7392 ( .IN1(g2081), .IN2(n2045), .IN3(n4474), .IN4(n3953), .Q(g20953) );
  OA22X1_S38584 U7393 ( .IN1(g2078), .IN2(n2045), .IN3(n4400), .IN4(n3953), .Q(g20934) );
  OA22X1_S38584 U7394 ( .IN1(g1411), .IN2(n1943), .IN3(n4417), .IN4(n3973), .Q(g20913) );
  OA22X1_S38584 U7395 ( .IN1(g1408), .IN2(n1943), .IN3(n4395), .IN4(n3973), .Q(g21070) );
  OA22X1_S38584 U7396 ( .IN1(g1405), .IN2(n1943), .IN3(n4475), .IN4(n3973), .Q(g21052) );
  OA22X1_S38584 U7397 ( .IN1(g1402), .IN2(n1943), .IN3(n4469), .IN4(n3973), .Q(g21033) );
  OA22X1_S38584 U7398 ( .IN1(g1399), .IN2(n1943), .IN3(n4411), .IN4(n3973), .Q(g21015) );
  OA22X1_S38584 U7399 ( .IN1(g1396), .IN2(n1943), .IN3(n4401), .IN4(n3973), .Q(g20993) );
  OA22X1_S38584 U7400 ( .IN1(g1393), .IN2(n1943), .IN3(n4412), .IN4(n3973), .Q(g20972) );
  OA22X1_S38584 U7401 ( .IN1(g1390), .IN2(n1943), .IN3(n4421), .IN4(n3973), .Q(g20949) );
  OA22X1_S38584 U7402 ( .IN1(g1387), .IN2(n1943), .IN3(n4476), .IN4(n3973), .Q(g20925) );
  OA22X1_S38584 U7403 ( .IN1(g1384), .IN2(n1943), .IN3(n4402), .IN4(n3973), .Q(g20910) );
  OA22X1_S38584 U7404 ( .IN1(g725), .IN2(n1842), .IN3(n4418), .IN4(n3993), .Q(g20894)
         );
  OA22X1_S38584 U7405 ( .IN1(g722), .IN2(n1842), .IN3(n4396), .IN4(n3993), .Q(g21051)
         );
  OA22X1_S38584 U7406 ( .IN1(g719), .IN2(n1842), .IN3(n4477), .IN4(n3993), .Q(g21031)
         );
  OA22X1_S38584 U7407 ( .IN1(g716), .IN2(n1842), .IN3(n4470), .IN4(n3993), .Q(g21009)
         );
  OA22X1_S38584 U7408 ( .IN1(g713), .IN2(n1842), .IN3(n4413), .IN4(n3993), .Q(g20989)
         );
  OA22X1_S38584 U7409 ( .IN1(g710), .IN2(n1842), .IN3(n4403), .IN4(n3993), .Q(g20966)
         );
  OA22X1_S38584 U7410 ( .IN1(g707), .IN2(n1842), .IN3(n4414), .IN4(n3993), .Q(g20944)
         );
  OA22X1_S38584 U7411 ( .IN1(g704), .IN2(n1842), .IN3(n4422), .IN4(n3993), .Q(g20921)
         );
  OA22X1_S38584 U7412 ( .IN1(g701), .IN2(n1842), .IN3(n4478), .IN4(n3993), .Q(g20901)
         );
  OA22X1_S38584 U7413 ( .IN1(g698), .IN2(n1842), .IN3(n4404), .IN4(n3993), .Q(g20891)
         );
  OA21X1 U7414 ( .IN1(g2812), .IN2(n4152), .IN3(n4153), .Q(g22269) );
  NOR2X0 U7415 ( .IN1(n4147), .IN2(n4306), .QN(n4152) );
  OA21X1 U7416 ( .IN1(g2118), .IN2(n4158), .IN3(n4159), .Q(g22249) );
  NOR2X0 U7417 ( .IN1(n4151), .IN2(n4307), .QN(n4158) );
  OA21X1 U7418 ( .IN1(g1424), .IN2(n4164), .IN3(n4165), .Q(g22234) );
  NOR2X0 U7419 ( .IN1(n4157), .IN2(n4308), .QN(n4164) );
  OA21X1 U7420 ( .IN1(g738), .IN2(n4167), .IN3(n4168), .Q(g22218) );
  NOR2X0 U7421 ( .IN1(n4163), .IN2(n4309), .QN(n4167) );
  OA22X1_S38584 U7422 ( .IN1(g2234), .IN2(n2086), .IN3(n4287), .IN4(n4170), .Q(g22154) );
  OA22X1_S38584 U7423 ( .IN1(g2233), .IN2(n2084), .IN3(n4287), .IN4(n4172), .Q(g22140) );
  OA22X1_S38584 U7424 ( .IN1(g2231), .IN2(n2086), .IN3(n4563), .IN4(n4170), .Q(g22139) );
  OA22X1_S38584 U7425 ( .IN1(g2230), .IN2(n2084), .IN3(n4563), .IN4(n4172), .Q(g22117) );
  OA22X1_S38584 U7426 ( .IN1(g2228), .IN2(n2086), .IN3(n4555), .IN4(n4170), .Q(g22116) );
  OA22X1_S38584 U7427 ( .IN1(g2227), .IN2(n2084), .IN3(n4555), .IN4(n4172), .Q(g22099) );
  OA22X1_S38584 U7428 ( .IN1(test_so74), .IN2(n2086), .IN3(n4325), .IN4(n4170), .Q(
        g22098) );
  OA22X1_S38584 U7429 ( .IN1(g2224), .IN2(n2084), .IN3(n4325), .IN4(n4172), .Q(g22078) );
  OA22X1_S38584 U7430 ( .IN1(g2222), .IN2(n2086), .IN3(n4389), .IN4(n4170), .Q(g22077) );
  OA22X1_S38584 U7431 ( .IN1(g2221), .IN2(n2084), .IN3(n4389), .IN4(n4172), .Q(g22061) );
  OA22X1_S38584 U7432 ( .IN1(g2219), .IN2(n2086), .IN3(n4319), .IN4(n4170), .Q(g22060) );
  OA22X1_S38584 U7433 ( .IN1(g2218), .IN2(n2084), .IN3(n4319), .IN4(n4172), .Q(g22045) );
  OA22X1_S38584 U7434 ( .IN1(g2210), .IN2(n2086), .IN3(n4373), .IN4(n4170), .Q(g22193) );
  OA22X1_S38584 U7435 ( .IN1(g2209), .IN2(n2084), .IN3(n4373), .IN4(n4172), .Q(g22183) );
  OA22X1_S38584 U7436 ( .IN1(g2207), .IN2(n2086), .IN3(n4377), .IN4(n4170), .Q(g22182) );
  OA22X1_S38584 U7437 ( .IN1(g2206), .IN2(n2084), .IN3(n4377), .IN4(n4172), .Q(g22170) );
  OA22X1_S38584 U7438 ( .IN1(g1540), .IN2(n1984), .IN3(n4288), .IN4(n4173), .Q(g22131) );
  OA22X1_S38584 U7439 ( .IN1(g1539), .IN2(n1982), .IN3(n4288), .IN4(n4175), .Q(g22114) );
  OA22X1_S38584 U7440 ( .IN1(test_so53), .IN2(n1984), .IN3(n4565), .IN4(n4173), .Q(
        g22113) );
  OA22X1_S38584 U7441 ( .IN1(g1536), .IN2(n1982), .IN3(n4565), .IN4(n4175), .Q(g22092) );
  OA22X1_S38584 U7442 ( .IN1(g1534), .IN2(n1984), .IN3(n4557), .IN4(n4173), .Q(g22091) );
  OA22X1_S38584 U7443 ( .IN1(g1533), .IN2(n1982), .IN3(n4557), .IN4(n4175), .Q(g22075) );
  OA22X1_S38584 U7444 ( .IN1(g1531), .IN2(n1984), .IN3(n4326), .IN4(n4173), .Q(g22074) );
  OA22X1_S38584 U7445 ( .IN1(g1530), .IN2(n1982), .IN3(n4326), .IN4(n4175), .Q(g22059) );
  OA22X1_S38584 U7446 ( .IN1(g1528), .IN2(n1984), .IN3(n4390), .IN4(n4173), .Q(g22058) );
  OA22X1_S38584 U7447 ( .IN1(g1527), .IN2(n1982), .IN3(n4390), .IN4(n4175), .Q(g22044) );
  OA22X1_S38584 U7448 ( .IN1(g1525), .IN2(n1984), .IN3(n4320), .IN4(n4173), .Q(g22043) );
  OA22X1_S38584 U7449 ( .IN1(g1524), .IN2(n1982), .IN3(n4320), .IN4(n4175), .Q(g22035) );
  OA22X1_S38584 U7450 ( .IN1(g1516), .IN2(n1984), .IN3(n4374), .IN4(n4173), .Q(g22179) );
  OA22X1_S38584 U7451 ( .IN1(test_so52), .IN2(n1982), .IN3(n4374), .IN4(n4175), .Q(
        g22167) );
  OA22X1_S38584 U7452 ( .IN1(g1513), .IN2(n1984), .IN3(n4378), .IN4(n4173), .Q(g22166) );
  OA22X1_S38584 U7453 ( .IN1(g1512), .IN2(n1982), .IN3(n4378), .IN4(n4175), .Q(g22149) );
  OA22X1_S38584 U7454 ( .IN1(g846), .IN2(n1882), .IN3(n4289), .IN4(n4176), .Q(g22105)
         );
  OA22X1_S38584 U7455 ( .IN1(g845), .IN2(n1880), .IN3(n4289), .IN4(n4178), .Q(g22089)
         );
  OA22X1_S38584 U7456 ( .IN1(g843), .IN2(n1882), .IN3(n4567), .IN4(n4176), .Q(g22088)
         );
  OA22X1_S38584 U7457 ( .IN1(g842), .IN2(n1880), .IN3(n4567), .IN4(n4178), .Q(g22068)
         );
  OA22X1_S38584 U7458 ( .IN1(g840), .IN2(n1882), .IN3(n4559), .IN4(n4176), .Q(g22067)
         );
  OA22X1_S38584 U7459 ( .IN1(test_so32), .IN2(n1880), .IN3(n4559), .IN4(n4178), .Q(
        g22056) );
  OA22X1_S38584 U7460 ( .IN1(g837), .IN2(n1882), .IN3(n4327), .IN4(n4176), .Q(g22055)
         );
  OA22X1_S38584 U7461 ( .IN1(g836), .IN2(n1880), .IN3(n4327), .IN4(n4178), .Q(g22042)
         );
  OA22X1_S38584 U7462 ( .IN1(g834), .IN2(n1882), .IN3(n4391), .IN4(n4176), .Q(g22041)
         );
  OA22X1_S38584 U7463 ( .IN1(g833), .IN2(n1880), .IN3(n4391), .IN4(n4178), .Q(g22034)
         );
  OA22X1_S38584 U7464 ( .IN1(g831), .IN2(n1882), .IN3(n4321), .IN4(n4176), .Q(g22033)
         );
  OA22X1_S38584 U7465 ( .IN1(g830), .IN2(n1880), .IN3(n4321), .IN4(n4178), .Q(g22029)
         );
  OA22X1_S38584 U7466 ( .IN1(g822), .IN2(n1882), .IN3(n4375), .IN4(n4176), .Q(g22163)
         );
  OA22X1_S38584 U7467 ( .IN1(g821), .IN2(n1880), .IN3(n4375), .IN4(n4178), .Q(g22146)
         );
  OA22X1_S38584 U7468 ( .IN1(g819), .IN2(n1882), .IN3(n4379), .IN4(n4176), .Q(g22145)
         );
  OA22X1_S38584 U7469 ( .IN1(g818), .IN2(n1880), .IN3(n4379), .IN4(n4178), .Q(g22126)
         );
  OA22X1_S38584 U7470 ( .IN1(g158), .IN2(n1778), .IN3(n4290), .IN4(n4179), .Q(g22080)
         );
  OA22X1_S38584 U7471 ( .IN1(g157), .IN2(n1776), .IN3(n4290), .IN4(n4180), .Q(g22065)
         );
  OA22X1_S38584 U7472 ( .IN1(g155), .IN2(n1778), .IN3(n4569), .IN4(n4179), .Q(g22064)
         );
  OA22X1_S38584 U7473 ( .IN1(g154), .IN2(n1776), .IN3(n4569), .IN4(n4180), .Q(g22049)
         );
  OA22X1_S38584 U7474 ( .IN1(g152), .IN2(n1778), .IN3(n4561), .IN4(n4179), .Q(g22048)
         );
  OA22X1_S38584 U7475 ( .IN1(g151), .IN2(n1776), .IN3(n4561), .IN4(n4180), .Q(g22039)
         );
  OA22X1_S38584 U7476 ( .IN1(g149), .IN2(n1778), .IN3(n4328), .IN4(n4179), .Q(g22038)
         );
  OA22X1_S38584 U7477 ( .IN1(g148), .IN2(n1776), .IN3(n4328), .IN4(n4180), .Q(g22032)
         );
  OA22X1_S38584 U7478 ( .IN1(g146), .IN2(n1778), .IN3(n4392), .IN4(n4179), .Q(g22031)
         );
  OA22X1_S38584 U7479 ( .IN1(g145), .IN2(n1776), .IN3(n4392), .IN4(n4180), .Q(g22028)
         );
  OA22X1_S38584 U7480 ( .IN1(g143), .IN2(n1778), .IN3(n4322), .IN4(n4179), .Q(g22027)
         );
  OA22X1_S38584 U7481 ( .IN1(g142), .IN2(n1776), .IN3(n4322), .IN4(n4180), .Q(g22025)
         );
  OA22X1_S38584 U7482 ( .IN1(g134), .IN2(n1778), .IN3(n4376), .IN4(n4179), .Q(g22142)
         );
  OA22X1_S38584 U7483 ( .IN1(g133), .IN2(n1776), .IN3(n4376), .IN4(n4180), .Q(g22123)
         );
  OA22X1_S38584 U7484 ( .IN1(g131), .IN2(n1778), .IN3(n4380), .IN4(n4179), .Q(g22122)
         );
  OA22X1_S38584 U7485 ( .IN1(g130), .IN2(n1776), .IN3(n4380), .IN4(n4180), .Q(g22100)
         );
  NBUFFX2 U7486 ( .IN(g2987), .Q(n4596) );
  OA21X1 U7487 ( .IN1(g2813), .IN2(n4148), .IN3(n3678), .Q(g22284) );
  NOR2X0 U7488 ( .IN1(n4147), .IN2(n4356), .QN(n4148) );
  OA21X1 U7489 ( .IN1(g2119), .IN2(n4154), .IN3(n3486), .Q(g22267) );
  NOR2X0 U7490 ( .IN1(n4151), .IN2(n4357), .QN(n4154) );
  OA21X1 U7491 ( .IN1(g1425), .IN2(n4160), .IN3(n3490), .Q(g22247) );
  NOR2X0 U7492 ( .IN1(n4157), .IN2(n4358), .QN(n4160) );
  OA21X1 U7493 ( .IN1(g739), .IN2(n4166), .IN3(n3494), .Q(g22231) );
  NOR2X0 U7494 ( .IN1(n4163), .IN2(n4359), .QN(n4166) );
  NOR2X0 U7495 ( .IN1(g3234), .IN2(DFF_1561_n1), .QN(g20884) );
  OA21X1 U7496 ( .IN1(test_so95), .IN2(n4145), .IN3(n4146), .Q(g22299) );
  NOR2X0 U7497 ( .IN1(n4147), .IN2(n4292), .QN(n4145) );
  OA21X1 U7498 ( .IN1(g2117), .IN2(n4149), .IN3(n4150), .Q(g22280) );
  NOR2X0 U7499 ( .IN1(n4151), .IN2(n4293), .QN(n4149) );
  OA21X1 U7500 ( .IN1(g1423), .IN2(n4155), .IN3(n4156), .Q(g22263) );
  NOR2X0 U7501 ( .IN1(n4157), .IN2(n4294), .QN(n4155) );
  OA21X1 U7502 ( .IN1(g737), .IN2(n4161), .IN3(n4162), .Q(g22242) );
  NOR2X0 U7503 ( .IN1(n4163), .IN2(n4295), .QN(n4161) );
  NOR2X0 U7504 ( .IN1(n4332), .IN2(g3231), .QN(n2419) );
  NBUFFX2 U7505 ( .IN(g3117), .Q(n4646) );
  NBUFFX2 U7506 ( .IN(g3129), .Q(g8106) );
  NBUFFX2 U7507 ( .IN(g3117), .Q(g8030) );
  NBUFFX2 U7508 ( .IN(g3109), .Q(n4644) );
  NBUFFX2 U7509 ( .IN(g2950), .Q(n4650) );
  NBUFFX2 U7510 ( .IN(g3129), .Q(n4648) );
  NOR2X0 U7511 ( .IN1(n2164), .IN2(n4062), .QN(g25197) );
  XOR2X1 U7512 ( .IN1(n3747), .IN2(g2734), .Q(n4062) );
  NOR2X0 U7513 ( .IN1(n2164), .IN2(n4126), .QN(g23348) );
  XOR2X1 U7514 ( .IN1(n4106), .IN2(g2727), .Q(n4126) );
  NOR2X0 U7515 ( .IN1(n2164), .IN2(n4217), .QN(g20789) );
  XOR2X1 U7516 ( .IN1(n4186), .IN2(g2714), .Q(n4217) );
  NOR2X0 U7517 ( .IN1(n2062), .IN2(n4063), .QN(g25194) );
  XOR2X1 U7518 ( .IN1(n3755), .IN2(g2040), .Q(n4063) );
  NOR2X0 U7519 ( .IN1(n2062), .IN2(n4127), .QN(g23339) );
  XOR2X1 U7520 ( .IN1(n4109), .IN2(g2033), .Q(n4127) );
  NOR2X0 U7521 ( .IN1(n2062), .IN2(n4218), .QN(g20752) );
  XOR2X1 U7522 ( .IN1(n4189), .IN2(g2020), .Q(n4218) );
  NOR2X0 U7523 ( .IN1(n1960), .IN2(n4067), .QN(g25189) );
  XOR2X1 U7524 ( .IN1(n3785), .IN2(g1346), .Q(n4067) );
  NOR2X0 U7525 ( .IN1(n1960), .IN2(n4131), .QN(g23329) );
  XOR2X1 U7526 ( .IN1(n4112), .IN2(g1339), .Q(n4131) );
  NOR2X0 U7527 ( .IN1(n1960), .IN2(n4219), .QN(g20717) );
  XOR2X1 U7528 ( .IN1(n4192), .IN2(g1326), .Q(n4219) );
  NOR2X0 U7529 ( .IN1(n1859), .IN2(n4068), .QN(g25185) );
  XOR2X1 U7530 ( .IN1(n3815), .IN2(g660), .Q(n4068) );
  NOR2X0 U7531 ( .IN1(n1859), .IN2(n4132), .QN(g23324) );
  XOR2X1 U7532 ( .IN1(n4115), .IN2(g653), .Q(n4132) );
  NOR2X0 U7533 ( .IN1(n1859), .IN2(n4220), .QN(g20682) );
  XOR2X1 U7534 ( .IN1(n4135), .IN2(g640), .Q(n4220) );
  OAI22X1 U7535 ( .IN1(n4299), .IN2(g2628), .IN3(n4352), .IN4(n4600), .QN(
        g18780) );
  OAI22X1 U7536 ( .IN1(n4366), .IN2(g1934), .IN3(n4311), .IN4(n4612), .QN(
        g18743) );
  OAI22X1 U7537 ( .IN1(n4300), .IN2(g1240), .IN3(n4353), .IN4(n4624), .QN(
        g18707) );
  OAI22X1 U7538 ( .IN1(n4313), .IN2(g554), .IN3(n4360), .IN4(n4634), .QN(
        g18678) );
  NAND2X0 U7539 ( .IN1(n1582), .IN2(DFF_1562_n1), .QN(n4263) );

  // Trigger ----------------------
  NOR2X0 Trojan1 ( .IN1(n3065), .IN2(n3016), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(n3023), .IN2(n3000), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(n3008), .IN2(n3068), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(n3128), .IN2(n3036), .QN(Tj_OUT4) );
  AND4X1 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT1), .IN3(Tj_OUT3), .IN4(Tj_OUT4), .Q(Tj_OUT1234) );

  NOR2X0 Trojan5 ( .IN1(n3758), .IN2(n3788), .QN(Tj_OUT5) );
  NOR2X0 Trojan6 ( .IN1(n3751), .IN2(n3749), .QN(Tj_OUT6) );
  NOR2X0 Trojan7 ( .IN1(n2792), .IN2(n2632), .QN(Tj_OUT7) );
  NOR2X0 Trojan8 ( .IN1(n2351), .IN2(n2430), .QN(Tj_OUT8) );
  AND4X1 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(Tj_OUT8), .Q(Tj_OUT5678) );

  AND2X1 Trojan_CLK_NOT ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .Q(Tj_Trigger) );

  // Payload ----------------------
  OR2X1 Trojan_Payload ( .IN1(Tj_Trigger), .IN2(n4263), .Q(n4263_Tj_Payload) );




endmodule

